// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.4.1.213
// Netlist written on Mon May  2 19:28:54 2016
//
// Verilog Description of module UniboardTop
//

module UniboardTop (uart_rx, uart_tx, status_led, clk_12MHz, Stepper_X_Step, 
            Stepper_X_Dir, Stepper_X_M0, Stepper_X_M1, Stepper_X_M2, 
            Stepper_X_En, Stepper_X_nFault, Stepper_Y_Step, Stepper_Y_Dir, 
            Stepper_Y_M0, Stepper_Y_M1, Stepper_Y_M2, Stepper_Y_En, 
            Stepper_Y_nFault, Stepper_Z_Step, Stepper_Z_Dir, Stepper_Z_M0, 
            Stepper_Z_M1, Stepper_Z_M2, Stepper_Z_En, Stepper_Z_nFault, 
            Stepper_A_Step, Stepper_A_Dir, Stepper_A_M0, Stepper_A_M1, 
            Stepper_A_M2, Stepper_A_En, Stepper_A_nFault, limit, expansion1, 
            expansion2, expansion3, expansion4, expansion5, signal_light, 
            encoder_ra, encoder_rb, encoder_ri, encoder_la, encoder_lb, 
            encoder_li, rc_ch1, rc_ch2, rc_ch3, rc_ch4, rc_ch7, 
            rc_ch8, motor_pwm_l, motor_pwm_r, xbee_pause, debug) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(362[8:19])
    input uart_rx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[13:20])
    output uart_tx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[14:21])
    output [2:0]status_led;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    input clk_12MHz;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    output Stepper_X_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(368[17:31])
    output Stepper_X_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:30])
    output Stepper_X_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:29])
    output Stepper_X_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    output Stepper_X_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    output Stepper_X_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    input Stepper_X_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[16:32])
    output Stepper_Y_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(376[17:31])
    output Stepper_Y_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:30])
    output Stepper_Y_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:29])
    output Stepper_Y_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    output Stepper_Y_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    output Stepper_Y_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    input Stepper_Y_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[16:32])
    output Stepper_Z_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(384[17:31])
    output Stepper_Z_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:30])
    output Stepper_Z_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:29])
    output Stepper_Z_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    output Stepper_Z_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    output Stepper_Z_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    input Stepper_Z_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[16:32])
    output Stepper_A_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(392[17:31])
    output Stepper_A_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:30])
    output Stepper_A_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:29])
    output Stepper_A_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    output Stepper_A_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    output Stepper_A_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    input Stepper_A_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[16:32])
    input [3:0]limit;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    output expansion1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[14:24])
    output expansion2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    output expansion3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    inout expansion4;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[13:23])
    input expansion5 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    output signal_light;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[14:26])
    input encoder_ra;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(408[13:23])
    input encoder_rb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    input encoder_ri;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    input encoder_la;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    input encoder_lb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    input encoder_li;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    input rc_ch1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(415[13:19])
    input rc_ch2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    input rc_ch3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    input rc_ch4;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    input rc_ch7;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    input rc_ch8;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    output motor_pwm_l;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(422[14:25])
    output motor_pwm_r;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    input xbee_pause;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[13:23])
    output [8:0]debug;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [127:0]select /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(455[15:21])
    wire n33384 /* synthesis nomerge= */ ;
    wire [15:0]battery_voltage;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(18[20:35])
    
    wire VCC_net, uart_rx_c, uart_tx_c, Stepper_X_Step_c, Stepper_X_Dir_c, 
        Stepper_X_M0_c_0, Stepper_X_M1_c_1, Stepper_X_M2_c_2, Stepper_X_En_c, 
        Stepper_X_nFault_c, Stepper_Y_Step_c, Stepper_Y_Dir_c, Stepper_Y_M0_c_0, 
        Stepper_Y_M1_c_1, Stepper_Y_M2_c_2, Stepper_Y_En_c, Stepper_Y_nFault_c, 
        Stepper_Z_Step_c, Stepper_Z_Dir_c, Stepper_Z_M0_c_0, Stepper_Z_M1_c_1, 
        Stepper_Z_M2_c_2, Stepper_Z_En_c, Stepper_Z_nFault_c, Stepper_A_Step_c, 
        Stepper_A_Dir_c, Stepper_A_M0_c_0, Stepper_A_M1_c_1, Stepper_A_M2_c_2, 
        Stepper_A_En_c, Stepper_A_nFault_c, limit_c_3, limit_c_2, limit_c_1, 
        limit_c_0, expansion1_c_9, expansion2_c_10, expansion3_c_11, 
        expansion5_c, signal_light_c, encoder_ra_c, encoder_rb_c, encoder_ri_c, 
        encoder_la_c, encoder_lb_c, encoder_li_c, rc_ch1_c, rc_ch2_c, 
        rc_ch3_c, rc_ch4_c, rc_ch7_c, rc_ch8_c, n11073, xbee_pause_c, 
        debug_c_7, debug_c_5, debug_c_4, debug_c_3, debug_c_2, debug_c_0;
    wire [31:0]databus;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(451[14:21])
    wire [2:0]reg_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(452[13:21])
    wire [7:0]register_addr;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    
    wire rw, n14454, n14547;
    wire [15:0]reset_count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(458[13:24])
    
    wire timeout_pause;
    wire [31:0]timeout_count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[13:26])
    
    wire prev_uart_rx, clk_255kHz, n27752, n27550, n14651, n1156, 
        n8, n9, n2;
    wire [31:0]n99_adj_1332;
    wire [7:0]n8635;
    
    wire n2_adj_605;
    wire [31:0]n100_adj_1351;
    wire [31:0]n658;
    
    wire n35;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    wire [31:0]databus_out;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(55[13:24])
    
    wire n21209, n13, n21212, n14, n21214, n6, n15087, n2967, 
        n21220, n21222;
    wire [31:0]n1474;
    
    wire n12, n29902, n29257, n14523, n31446, n29827, n5834, n8507, 
        n9369, n2876, n2870, n14514, n14513, n3, n2_adj_606, n27445;
    wire [31:0]n5974;
    
    wire n29944, n2861, n2858, n10, n32, n13316, n3_adj_607, n8_adj_608, 
        n24, n2_adj_609, n9538, n4007, force_pause;
    wire [31:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(24[14:22])
    wire [31:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(24[14:22])
    
    wire clk_1Hz, prev_clk_1Hz;
    wire [31:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(31[13:23])
    wire [2:0]read_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(32[12:21])
    
    wire n46, n22396, n22390, n14146, n31410;
    wire [7:0]\register[0]_adj_971 ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    wire [7:0]read_value_adj_972;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(92[12:22])
    
    wire n22;
    wire [2:0]read_size_adj_973;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(93[12:21])
    
    wire n64, n32_adj_619, n16843, n16842, n34, n27536, n29237, 
        n3_adj_620, n27442, n2847, n14500, n16841, n241, n27428, 
        n9331;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire limit_latched, prev_limit_latched, step_clk, prev_step_clk;
    wire [31:0]read_value_adj_979;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_980;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select, n52, n17, n16, n15, n303, n31445, n31444, 
        n73, n18, n16013, n4181;
    wire [7:0]control_reg_adj_988;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]div_factor_reg_adj_989;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg_adj_990;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire limit_latched_adj_656, prev_limit_latched_adj_657, int_step, 
        step_clk_adj_658, prev_step_clk_adj_659;
    wire [31:0]read_value_adj_991;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_992;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_694, n4, n52_adj_695;
    wire [31:0]n224_adj_995;
    
    wire n27169, n27168, n27167, n27166, n8402, n31443, n27165;
    wire [31:0]n4095;
    
    wire n27164, n27163, n8_adj_697, n8368, n14_adj_698, n13_adj_699, 
        n27162, n27161, n2_adj_700, n33388, n27160, n27159, n3_adj_701;
    wire [31:0]steps_reg_adj_1029;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire limit_latched_adj_702, prev_limit_latched_adj_703;
    wire [31:0]read_value_adj_1030;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_1031;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_738, n8_adj_739, n11, n8_adj_740, n2_adj_741, 
        n13957, n9305, n13948, n2_adj_742, n8056, n13941, n33387;
    wire [31:0]n580_adj_1049;
    
    wire n13939, n9301, n5;
    wire [7:0]control_reg_adj_1066;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire limit_latched_adj_744, prev_limit_latched_adj_745;
    wire [31:0]read_value_adj_1069;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_1070;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_780, n29838;
    wire [31:0]n224_adj_1073;
    
    wire n8298, n8_adj_813, n31411, n8_adj_814, n8_adj_815;
    wire [31:0]n3922;
    
    wire n27543, n13917, n2_adj_816, n9484, n29784, n9297, n29492, 
        n13908, n2_adj_817, n8264, n8_adj_818, n31409, n2824;
    wire [31:0]\register[1]_adj_1105 ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(58[14:22])
    
    wire qreset;
    wire [31:0]read_value_adj_1107;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(65[13:23])
    wire [2:0]read_size_adj_1108;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(66[12:21])
    
    wire prev_select_adj_853;
    wire [31:0]read_value_adj_1115;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(65[13:23])
    wire [2:0]read_size_adj_1116;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(66[12:21])
    
    wire prev_select_adj_888;
    wire [7:0]\register[1]_adj_1129 ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(17[12:20])
    wire [7:0]\register[0]_adj_1130 ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(17[12:20])
    wire [7:0]read_value_adj_1131;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(26[12:22])
    wire [2:0]read_size_adj_1132;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(27[12:21])
    
    wire prev_select_adj_898, n176, n31413, n13834, n29235, n29294, 
        n29301, n9_adj_899, n29293, n2_adj_900, n3_adj_901, n2_adj_902, 
        n2_adj_903, n8_adj_904;
    wire [14:0]n33692;
    
    wire n8_adj_906, n12211, n31412, n31436, n31435, n31432, n31428, 
        n31427, n31426, n31425, n6_adj_907, n33385, n27680, n29818, 
        n1, n2_adj_908, n8_adj_909, n14_adj_910, n2_adj_911, n2_adj_912, 
        n8_adj_913, n24146, n29792, n2_adj_914, n29847, n2_adj_915, 
        n8_adj_916, n2_adj_917, n2_adj_918, n8_adj_919, n8_adj_920, 
        n29811, n2_adj_921, n8_adj_922, n2_adj_923, n8_adj_924, n29789, 
        n2_adj_925, n2_adj_926, n12149, n8_adj_927, n8_adj_928, n2_adj_929, 
        n2_adj_930, n8_adj_931, n3_adj_932, n2_adj_933, n2_adj_934, 
        n8_adj_935, n29170, n2_adj_936, n29530, n26435, n29840;
    wire [7:0]n8653;
    
    wire n56, n26434, n66, n2_adj_937, n22484, n9_adj_938, n8194, 
        n26433, n14783, n31601, n27541, n11236;
    wire [31:0]n6779;
    
    wire n30, n26432, n26431, n31596, n17035, select_clk, n9379, 
        n26430, n31591, n31590, n26429, n26428, n26427, n31588, 
        n31422, n26426;
    wire [1:0]n33625;
    
    wire n31582, n42, n40, n38, n36, n34_adj_940, expansion4_out, 
        n31576, n30_adj_941, n29, n30306, n26, n29271, n31571, 
        n26425, n29137, n31556, n11008, n33386, n11209, n2_adj_942, 
        n2_adj_943, n29264, n6_adj_944, n12369, n31541, n31540, 
        n29334, n31537, n7917, n21503, n31533, n27564;
    wire [2:0]quadA_delayed_adj_1219;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    wire [2:0]quadB_delayed_adj_1220;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    
    wire n31530, n8160, n33390, n27753, n8_adj_945, n8_adj_946, 
        n29114, n11007, n31526, n12159, n9581, n9548, n9542, n3_adj_947, 
        n30304, n31512, n7882, n29200, n29067, n28827, n29057, 
        n29054, n29066, n29064, n29051, n29053, n29055, n31504, 
        n29068, n29058, n31502, n27547, n29069, n29072, n31501, 
        n29071, n27465, n31497, n29059, n29060, n29065, n29061, 
        n29063, n31407, n29056, n29052, n31408, n29050, n29062, 
        n29049, n29070, n29295, n29221, n3_adj_948, n31421, n29832, 
        n7847, n27484, n8090, n29258, n31483, n29113, n27250, 
        n31478, n31477, n31474, n31473, n31420, n31471, n31470, 
        n31466, n16765, n31465, n29332, n31464, n31419, n31463, 
        n26424, n26423, n26422, n26421, n31457, n26420, n107;
    wire [3:0]state_adj_1308;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n29048, n26890, n26889, n13156, n27785, n31450, n26888, 
        n26887, n29830, n26886, n26885, n31449, n26884, n16764, 
        n31447, n29786;
    
    VHI i2 (.Z(VCC_net));
    ExpansionGPIO gpio (.read_value({read_value_adj_1131}), .debug_c_c(debug_c_c), 
            .n2870(n2870), .n29221(n29221), .n13948(n13948), .n31512(n31512), 
            .\databus[0] (databus[0]), .\read_size[0] (read_size_adj_1132[0]), 
            .n27680(n27680), .prev_select(prev_select_adj_898), .\select[5] (select[5]), 
            .expansion1_c_9(expansion1_c_9), .n31436(n31436), .n56(n56), 
            .expansion2_c_10(expansion2_c_10), .expansion3_c_11(expansion3_c_11), 
            .\databus[1] (databus[1]), .\databus[2] (databus[2]), .\databus[3] (databus[3]), 
            .\register[0][4] (\register[0]_adj_1130 [4]), .\databus[4] (databus[4]), 
            .\register[0][5] (\register[0]_adj_1130 [5]), .\databus[5] (databus[5]), 
            .\databus[6] (databus[6]), .\databus[7] (databus[7]), .n16013(n16013), 
            .\register[1][4] (\register[1]_adj_1129 [4]), .\register[1][5] (\register[1]_adj_1129 [5]), 
            .n12369(n12369), .n31407(n31407), .\register_addr[0] (register_addr[0]), 
            .n24146(n24146), .n11008(n11008), .n11007(n11007)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(694[18] 705[38])
    IFS1P3DX prev_uart_rx_58 (.D(uart_rx_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(battery_voltage[15]), .Q(prev_uart_rx));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam prev_uart_rx_58.GSR = "ENABLED";
    FD1S3AX timeout_pause_60 (.D(n27785), .CK(debug_c_c), .Q(timeout_pause));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_pause_60.GSR = "ENABLED";
    LUT4 i1044_2_lut_rep_266_3_lut (.A(n22484), .B(reset_count[14]), .C(n8368), 
         .Z(n31410)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1044_2_lut_rep_266_3_lut.init = 16'hf7f7;
    LUT4 i15032_2_lut_2_lut_3_lut (.A(n22484), .B(reset_count[14]), .C(databus[4]), 
         .Z(n580_adj_1049[4])) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15032_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i2_3_lut_rep_269_4_lut (.A(n22484), .B(reset_count[14]), .C(n8507), 
         .D(select_clk), .Z(n31413)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_269_4_lut.init = 16'h0080;
    CCU2D add_31_9 (.A0(timeout_count[7]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[8]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26423), 
          .COUT(n26424), .S0(n658[7]), .S1(n658[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_9.INIT0 = 16'h5aaa;
    defparam add_31_9.INIT1 = 16'h5aaa;
    defparam add_31_9.INJECT1_0 = "NO";
    defparam add_31_9.INJECT1_1 = "NO";
    CCU2D add_31_7 (.A0(timeout_count[5]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[6]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26422), 
          .COUT(n26423), .S0(n658[5]), .S1(n658[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_7.INIT0 = 16'h5aaa;
    defparam add_31_7.INIT1 = 16'h5aaa;
    defparam add_31_7.INJECT1_0 = "NO";
    defparam add_31_7.INJECT1_1 = "NO";
    LUT4 i10292_2_lut_3_lut_4_lut (.A(n22484), .B(reset_count[14]), .C(n8090), 
         .D(n8056), .Z(n17035)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i10292_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i14815_2_lut_2_lut_3_lut (.A(n22484), .B(reset_count[14]), .C(n7882), 
         .Z(n241)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i14815_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i5445_3_lut_4_lut (.A(n22484), .B(reset_count[14]), .C(limit_latched_adj_744), 
         .D(prev_limit_latched_adj_745), .Z(n12211)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i5445_3_lut_4_lut.init = 16'h77f7;
    LUT4 i22482_3_lut_4_lut (.A(n22484), .B(reset_count[14]), .C(n73), 
         .D(state_adj_1308[2]), .Z(n14783)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i22482_3_lut_4_lut.init = 16'hff7f;
    LUT4 i22345_4_lut (.A(n29334), .B(reset_count[14]), .C(n13316), .D(n21503), 
         .Z(n30)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam i22345_4_lut.init = 16'h373f;
    LUT4 i1_2_lut_3_lut (.A(n22484), .B(reset_count[14]), .C(n9305), .Z(n14547)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_4_lut (.A(n22396), .B(n29332), .C(reset_count[6]), .D(reset_count[5]), 
         .Z(n29334)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(461[7:30])
    defparam i1_4_lut.init = 16'hfcec;
    LUT4 i1_3_lut_4_lut (.A(n22484), .B(reset_count[14]), .C(prev_limit_latched_adj_703), 
         .D(limit_latched_adj_702), .Z(n11209)) /* synthesis lut_function=(!(A (B (C+!(D))))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h7f77;
    LUT4 i15653_4_lut (.A(reset_count[0]), .B(reset_count[4]), .C(n6_adj_907), 
         .D(reset_count[3]), .Z(n22396)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i15653_4_lut.init = 16'hccc8;
    LUT4 i2_2_lut (.A(reset_count[1]), .B(reset_count[2]), .Z(n6_adj_907)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut (.A(reset_count[11]), .B(reset_count[12]), .C(reset_count[13]), 
         .Z(n13316)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(461[7:30])
    defparam i2_3_lut.init = 16'hfefe;
    VLO i1 (.Z(battery_voltage[15]));
    LUT4 i4_2_lut_3_lut (.A(n22484), .B(reset_count[14]), .C(debug_c_0), 
         .Z(qreset)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i4_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_3_lut_4_lut_adj_509 (.A(n22484), .B(reset_count[14]), .C(prev_limit_latched), 
         .D(limit_latched), .Z(n12159)) /* synthesis lut_function=(!(A (B (C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_509.init = 16'h7f77;
    LUT4 i5384_3_lut_4_lut (.A(n22484), .B(reset_count[14]), .C(limit_latched_adj_656), 
         .D(prev_limit_latched_adj_657), .Z(n12149)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i5384_3_lut_4_lut.init = 16'h77f7;
    LUT4 i22328_2_lut_3_lut (.A(n22484), .B(reset_count[14]), .C(n29786), 
         .Z(n2967)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i22328_2_lut_3_lut.init = 16'hf7f7;
    FD1P3IX timeout_count__i0 (.D(n100_adj_1351[0]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i0.GSR = "ENABLED";
    LUT4 i22331_2_lut_3_lut (.A(n22484), .B(reset_count[14]), .C(n29789), 
         .Z(n2876)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i22331_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i22334_2_lut_3_lut (.A(n22484), .B(reset_count[14]), .C(n29792), 
         .Z(n2861)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i22334_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i974_2_lut_3_lut (.A(n22484), .B(reset_count[14]), .C(n7917), 
         .Z(n2824)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i974_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1032_2_lut_rep_265_3_lut (.A(n22484), .B(reset_count[14]), .C(n8056), 
         .Z(n31409)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1032_2_lut_rep_265_3_lut.init = 16'hf7f7;
    LUT4 i10069_2_lut_3_lut_4_lut (.A(n22484), .B(reset_count[14]), .C(n8194), 
         .D(n8160), .Z(n16841)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i10069_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i1036_2_lut_rep_264_3_lut (.A(n22484), .B(reset_count[14]), .C(n8160), 
         .Z(n31408)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1036_2_lut_rep_264_3_lut.init = 16'hf7f7;
    CCU2D add_31_5 (.A0(timeout_count[3]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[4]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26421), 
          .COUT(n26422), .S0(n100_adj_1351[3]), .S1(n658[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_5.INIT0 = 16'h5aaa;
    defparam add_31_5.INIT1 = 16'h5aaa;
    defparam add_31_5.INJECT1_0 = "NO";
    defparam add_31_5.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_268_4_lut (.A(n22484), .B(reset_count[14]), .C(n7882), 
         .D(clk_255kHz), .Z(n31412)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_268_4_lut.init = 16'h0080;
    LUT4 i1_3_lut_rep_319_4_lut (.A(n22484), .B(reset_count[14]), .C(state_adj_1308[3]), 
         .D(state_adj_1308[2]), .Z(n31463)) /* synthesis lut_function=(!(((C (D))+!B)+!A)) */ ;
    defparam i1_3_lut_rep_319_4_lut.init = 16'h0888;
    LUT4 i2759_3_lut_4_lut (.A(n22484), .B(reset_count[14]), .C(prev_clk_1Hz), 
         .D(clk_1Hz), .Z(n9484)) /* synthesis lut_function=(!(A (B (C+!(D))))) */ ;
    defparam i2759_3_lut_4_lut.init = 16'h7f77;
    LUT4 i10070_2_lut_3_lut_4_lut (.A(n22484), .B(reset_count[14]), .C(n8298), 
         .D(n8264), .Z(n16842)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i10070_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i1040_2_lut_rep_267_3_lut (.A(n22484), .B(reset_count[14]), .C(n8264), 
         .Z(n31411)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1040_2_lut_rep_267_3_lut.init = 16'hf7f7;
    LUT4 i15230_2_lut_2_lut_3_lut (.A(n22484), .B(reset_count[14]), .C(n8507), 
         .Z(n107)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15230_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i10071_2_lut_3_lut_4_lut (.A(n22484), .B(reset_count[14]), .C(n8402), 
         .D(n8368), .Z(n16843)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i10071_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i14851_2_lut_2_lut_3_lut (.A(n22484), .B(reset_count[14]), .C(databus[2]), 
         .Z(n580_adj_1049[2])) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i14851_2_lut_2_lut_3_lut.init = 16'h8080;
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i2_3_lut_rep_288_4_lut (.A(select[3]), .B(n31502), .C(n31526), 
         .D(prev_select_adj_888), .Z(n31432)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam i2_3_lut_rep_288_4_lut.init = 16'h0080;
    LUT4 Select_4296_i10_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1115[1]), 
         .D(n33385), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4296_i10_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_3_lut_3_lut (.A(n31501), .B(n1474[17]), .C(n1474[20]), .Z(n27465)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i2_3_lut_3_lut.init = 16'hfdfd;
    LUT4 i22363_4_lut_4_lut (.A(n31501), .B(n4), .C(n5834), .D(n1474[14]), 
         .Z(n13834)) /* synthesis lut_function=(!((B (C+!(D))+!B !(D))+!A)) */ ;
    defparam i22363_4_lut_4_lut.init = 16'h2a00;
    LUT4 i2_3_lut_rep_469 (.A(n22484), .B(reset_count[14]), .C(n7882), 
         .D(clk_255kHz), .Z(n33388)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_469.init = 16'h0080;
    CCU2D add_19623_24 (.A0(timeout_count[31]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(battery_voltage[15]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27169), .S1(n7847));
    defparam add_19623_24.INIT0 = 16'h5555;
    defparam add_19623_24.INIT1 = 16'h0000;
    defparam add_19623_24.INJECT1_0 = "NO";
    defparam add_19623_24.INJECT1_1 = "NO";
    CCU2D add_19623_22 (.A0(timeout_count[29]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[30]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27168), .COUT(n27169));
    defparam add_19623_22.INIT0 = 16'h5555;
    defparam add_19623_22.INIT1 = 16'h5555;
    defparam add_19623_22.INJECT1_0 = "NO";
    defparam add_19623_22.INJECT1_1 = "NO";
    CCU2D add_19623_20 (.A0(timeout_count[27]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[28]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27167), .COUT(n27168));
    defparam add_19623_20.INIT0 = 16'h5555;
    defparam add_19623_20.INIT1 = 16'h5555;
    defparam add_19623_20.INJECT1_0 = "NO";
    defparam add_19623_20.INJECT1_1 = "NO";
    CCU2D add_19623_18 (.A0(timeout_count[25]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[26]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27166), .COUT(n27167));
    defparam add_19623_18.INIT0 = 16'h5aaa;
    defparam add_19623_18.INIT1 = 16'h5555;
    defparam add_19623_18.INJECT1_0 = "NO";
    defparam add_19623_18.INJECT1_1 = "NO";
    CCU2D add_19623_16 (.A0(timeout_count[23]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[24]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27165), .COUT(n27166));
    defparam add_19623_16.INIT0 = 16'h5aaa;
    defparam add_19623_16.INIT1 = 16'h5aaa;
    defparam add_19623_16.INJECT1_0 = "NO";
    defparam add_19623_16.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n31512), .B(prev_select_adj_780), 
         .C(n31466), .D(register_addr[5]), .Z(n2858)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h1000;
    CCU2D add_19623_14 (.A0(timeout_count[21]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[22]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27164), .COUT(n27165));
    defparam add_19623_14.INIT0 = 16'h5555;
    defparam add_19623_14.INIT1 = 16'h5555;
    defparam add_19623_14.INJECT1_0 = "NO";
    defparam add_19623_14.INJECT1_1 = "NO";
    CCU2D add_19623_12 (.A0(timeout_count[19]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[20]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27163), .COUT(n27164));
    defparam add_19623_12.INIT0 = 16'h5555;
    defparam add_19623_12.INIT1 = 16'h5aaa;
    defparam add_19623_12.INJECT1_0 = "NO";
    defparam add_19623_12.INJECT1_1 = "NO";
    CCU2D add_19623_10 (.A0(timeout_count[17]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[18]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27162), .COUT(n27163));
    defparam add_19623_10.INIT0 = 16'h5aaa;
    defparam add_19623_10.INIT1 = 16'h5555;
    defparam add_19623_10.INJECT1_0 = "NO";
    defparam add_19623_10.INJECT1_1 = "NO";
    CCU2D add_19623_8 (.A0(timeout_count[15]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[16]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27161), .COUT(n27162));
    defparam add_19623_8.INIT0 = 16'h5aaa;
    defparam add_19623_8.INIT1 = 16'h5aaa;
    defparam add_19623_8.INJECT1_0 = "NO";
    defparam add_19623_8.INJECT1_1 = "NO";
    CCU2D add_19623_6 (.A0(timeout_count[13]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[14]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27160), .COUT(n27161));
    defparam add_19623_6.INIT0 = 16'h5555;
    defparam add_19623_6.INIT1 = 16'h5555;
    defparam add_19623_6.INJECT1_0 = "NO";
    defparam add_19623_6.INJECT1_1 = "NO";
    CCU2D add_19623_4 (.A0(timeout_count[11]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[12]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27159), .COUT(n27160));
    defparam add_19623_4.INIT0 = 16'h5555;
    defparam add_19623_4.INIT1 = 16'h5555;
    defparam add_19623_4.INJECT1_0 = "NO";
    defparam add_19623_4.INJECT1_1 = "NO";
    LUT4 i22443_4_lut (.A(n29902), .B(n17), .C(n15), .D(n16), .Z(n27785)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i22443_4_lut.init = 16'h8000;
    CCU2D add_19623_2 (.A0(timeout_count[9]), .B0(timeout_count[8]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[10]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .COUT(n27159));
    defparam add_19623_2.INIT0 = 16'h7000;
    defparam add_19623_2.INIT1 = 16'h5aaa;
    defparam add_19623_2.INJECT1_0 = "NO";
    defparam add_19623_2.INJECT1_1 = "NO";
    LUT4 i22442_4_lut (.A(n29), .B(n42), .C(n38), .D(n30_adj_941), .Z(n29902)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i22442_4_lut.init = 16'h0001;
    LUT4 i7_4_lut (.A(timeout_count[16]), .B(timeout_count[25]), .C(timeout_count[15]), 
         .D(timeout_count[24]), .Z(n17)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i5_2_lut (.A(timeout_count[8]), .B(timeout_count[20]), .Z(n15)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5_2_lut.init = 16'h8888;
    LUT4 i6_4_lut (.A(timeout_count[17]), .B(timeout_count[9]), .C(timeout_count[23]), 
         .D(timeout_count[10]), .Z(n16)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i7_2_lut (.A(timeout_count[5]), .B(timeout_count[18]), .Z(n29)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(timeout_count[12]), .B(n40), .C(n34_adj_940), .D(timeout_count[19]), 
         .Z(n42)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(timeout_count[31]), .B(timeout_count[22]), .C(timeout_count[21]), 
         .D(timeout_count[28]), .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i16_4_lut.init = 16'hfffe;
    FD1P3AX reset_count_2669_2670__i1 (.D(n33692[0]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670__i1.GSR = "ENABLED";
    LUT4 i8_2_lut (.A(timeout_count[1]), .B(timeout_count[4]), .Z(n30_adj_941)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i18_4_lut (.A(timeout_count[6]), .B(n36), .C(n26), .D(timeout_count[2]), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i12_4_lut (.A(timeout_count[14]), .B(timeout_count[11]), .C(timeout_count[30]), 
         .D(timeout_count[13]), .Z(n34_adj_940)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(timeout_count[29]), .B(timeout_count[26]), .C(timeout_count[7]), 
         .D(timeout_count[3]), .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(timeout_count[0]), .B(timeout_count[27]), .Z(n26)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_rep_357 (.A(reset_count[14]), .B(reset_count[12]), .C(reset_count[13]), 
         .D(n29264), .Z(n31501)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam i1_4_lut_rep_357.init = 16'hfaea;
    LUT4 i15746_1_lut_rep_329_4_lut (.A(reset_count[14]), .B(reset_count[12]), 
         .C(reset_count[13]), .D(n29264), .Z(n31473)) /* synthesis lut_function=(!(A+(B (C)+!B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam i15746_1_lut_rep_329_4_lut.init = 16'h0515;
    LUT4 i15_2_lut_rep_300_3_lut_4_lut (.A(register_addr[4]), .B(n31533), 
         .C(rw), .D(select[3]), .Z(n31444)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam i15_2_lut_rep_300_3_lut_4_lut.init = 16'hd000;
    LUT4 i114_2_lut_3_lut_4_lut (.A(register_addr[4]), .B(n31533), .C(prev_select_adj_853), 
         .D(select[3]), .Z(n14146)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam i114_2_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 Select_4301_i6_2_lut_3_lut_4_lut (.A(register_addr[4]), .B(n31533), 
         .C(read_size_adj_1108[2]), .D(select[3]), .Z(n6)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4301_i6_2_lut_3_lut_4_lut.init = 16'hd000;
    LUT4 i15_2_lut_rep_303_3_lut_4_lut (.A(register_addr[4]), .B(n31533), 
         .C(rw), .D(select[3]), .Z(n31447)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam i15_2_lut_rep_303_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4308_i9_2_lut_3_lut_4_lut (.A(register_addr[4]), .B(n31533), 
         .C(read_size_adj_1116[0]), .D(select[3]), .Z(n9)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4308_i9_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i114_2_lut_3_lut_4_lut_adj_510 (.A(register_addr[4]), .B(n31533), 
         .C(prev_select_adj_888), .D(select[3]), .Z(n15087)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam i114_2_lut_3_lut_4_lut_adj_510.init = 16'h0200;
    LUT4 i2_3_lut_rep_467 (.A(n22484), .B(reset_count[14]), .C(n7882), 
         .D(clk_255kHz), .Z(n33386)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_467.init = 16'h0080;
    LUT4 i2_3_lut_rep_468 (.A(n22484), .B(reset_count[14]), .C(n7882), 
         .D(clk_255kHz), .Z(n33387)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_468.init = 16'h0080;
    LUT4 i22421_2_lut_rep_368 (.A(n22484), .B(reset_count[14]), .Z(n31512)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i22421_2_lut_rep_368.init = 16'h7777;
    CCU2D add_31_3 (.A0(timeout_count[1]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[2]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26420), 
          .COUT(n26421), .S0(n100_adj_1351[1]), .S1(n100_adj_1351[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_3.INIT0 = 16'h5aaa;
    defparam add_31_3.INIT1 = 16'h5aaa;
    defparam add_31_3.INJECT1_0 = "NO";
    defparam add_31_3.INJECT1_1 = "NO";
    LUT4 Select_4232_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[27]), 
         .D(n33385), .Z(n8_adj_814)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4232_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    CCU2D add_31_1 (.A0(battery_voltage[15]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[0]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .COUT(n26420), .S1(n100_adj_1351[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_1.INIT0 = 16'hF000;
    defparam add_31_1.INIT1 = 16'h5555;
    defparam add_31_1.INJECT1_0 = "NO";
    defparam add_31_1.INJECT1_1 = "NO";
    LUT4 i14774_2_lut (.A(reset_count[9]), .B(reset_count[10]), .Z(n21503)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14774_2_lut.init = 16'h8888;
    IB xbee_pause_pad (.I(xbee_pause), .O(xbee_pause_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[13:23])
    IB rc_ch8_pad (.I(rc_ch8), .O(rc_ch8_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    IB rc_ch7_pad (.I(rc_ch7), .O(rc_ch7_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    IB rc_ch4_pad (.I(rc_ch4), .O(rc_ch4_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    IB rc_ch3_pad (.I(rc_ch3), .O(rc_ch3_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    IB rc_ch2_pad (.I(rc_ch2), .O(rc_ch2_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    IB rc_ch1_pad (.I(rc_ch1), .O(rc_ch1_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(415[13:19])
    IB encoder_li_pad (.I(encoder_li), .O(encoder_li_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    IB encoder_lb_pad (.I(encoder_lb), .O(encoder_lb_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    IB encoder_la_pad (.I(encoder_la), .O(encoder_la_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    IB encoder_ri_pad (.I(encoder_ri), .O(encoder_ri_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    IB encoder_rb_pad (.I(encoder_rb), .O(encoder_rb_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    IB encoder_ra_pad (.I(encoder_ra), .O(encoder_ra_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(408[13:23])
    IB expansion5_pad (.I(expansion5), .O(expansion5_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    IB limit_pad_0 (.I(limit[0]), .O(limit_c_0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB limit_pad_1 (.I(limit[1]), .O(limit_c_1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB limit_pad_2 (.I(limit[2]), .O(limit_c_2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB limit_pad_3 (.I(limit[3]), .O(limit_c_3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB Stepper_A_nFault_pad (.I(Stepper_A_nFault), .O(Stepper_A_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[16:32])
    IB Stepper_Z_nFault_pad (.I(Stepper_Z_nFault), .O(Stepper_Z_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[16:32])
    IB Stepper_Y_nFault_pad (.I(Stepper_Y_nFault), .O(Stepper_Y_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[16:32])
    IB Stepper_X_nFault_pad (.I(Stepper_X_nFault), .O(Stepper_X_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[16:32])
    IB debug_c_pad (.I(clk_12MHz), .O(debug_c_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    IB uart_rx_pad (.I(uart_rx), .O(uart_rx_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[13:20])
    OB debug_pad_0 (.I(debug_c_0), .O(debug[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_1 (.I(n11073), .O(debug[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_2 (.I(debug_c_2), .O(debug[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_3 (.I(debug_c_3), .O(debug[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_4 (.I(debug_c_4), .O(debug[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_5 (.I(debug_c_5), .O(debug[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_6 (.I(n31512), .O(debug[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_7 (.I(debug_c_7), .O(debug[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_8 (.I(debug_c_c), .O(debug[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB motor_pwm_r_pad (.I(n11073), .O(motor_pwm_r));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    OB motor_pwm_l_pad (.I(n11073), .O(motor_pwm_l));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(422[14:25])
    OB signal_light_pad (.I(signal_light_c), .O(signal_light));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[14:26])
    OB expansion3_pad (.I(expansion3_c_11), .O(expansion3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    OB expansion2_pad (.I(expansion2_c_10), .O(expansion2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    OB expansion1_pad (.I(expansion1_c_9), .O(expansion1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[14:24])
    OB Stepper_A_En_pad (.I(Stepper_A_En_c), .O(Stepper_A_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    OB Stepper_A_M2_pad (.I(Stepper_A_M2_c_2), .O(Stepper_A_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    OB Stepper_A_M1_pad (.I(Stepper_A_M1_c_1), .O(Stepper_A_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    OB Stepper_A_M0_pad (.I(Stepper_A_M0_c_0), .O(Stepper_A_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:29])
    OB Stepper_A_Dir_pad (.I(Stepper_A_Dir_c), .O(Stepper_A_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:30])
    OB Stepper_A_Step_pad (.I(Stepper_A_Step_c), .O(Stepper_A_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(392[17:31])
    OB Stepper_Z_En_pad (.I(Stepper_Z_En_c), .O(Stepper_Z_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    OB Stepper_Z_M2_pad (.I(Stepper_Z_M2_c_2), .O(Stepper_Z_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    OB Stepper_Z_M1_pad (.I(Stepper_Z_M1_c_1), .O(Stepper_Z_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    OB Stepper_Z_M0_pad (.I(Stepper_Z_M0_c_0), .O(Stepper_Z_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:29])
    OB Stepper_Z_Dir_pad (.I(Stepper_Z_Dir_c), .O(Stepper_Z_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:30])
    CCU2D add_31_33 (.A0(timeout_count[31]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(battery_voltage[15]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26435), 
          .S0(n658[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_33.INIT0 = 16'h5aaa;
    defparam add_31_33.INIT1 = 16'h0000;
    defparam add_31_33.INJECT1_0 = "NO";
    defparam add_31_33.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut_4_lut (.A(n31512), .B(n31582), .C(n31477), .D(register_addr[1]), 
         .Z(n9542)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i2_3_lut_4_lut_4_lut.init = 16'h4440;
    LUT4 Select_4235_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[26]), 
         .D(n33385), .Z(n8_adj_913)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4235_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    OB Stepper_Z_Step_pad (.I(Stepper_Z_Step_c), .O(Stepper_Z_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(384[17:31])
    OB Stepper_Y_En_pad (.I(Stepper_Y_En_c), .O(Stepper_Y_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    CCU2D add_31_31 (.A0(timeout_count[29]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[30]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26434), 
          .COUT(n26435), .S0(n658[29]), .S1(n658[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_31.INIT0 = 16'h5aaa;
    defparam add_31_31.INIT1 = 16'h5aaa;
    defparam add_31_31.INJECT1_0 = "NO";
    defparam add_31_31.INJECT1_1 = "NO";
    CCU2D add_31_17 (.A0(timeout_count[15]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[16]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26427), 
          .COUT(n26428), .S0(n658[15]), .S1(n658[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_17.INIT0 = 16'h5aaa;
    defparam add_31_17.INIT1 = 16'h5aaa;
    defparam add_31_17.INJECT1_0 = "NO";
    defparam add_31_17.INJECT1_1 = "NO";
    CCU2D add_31_29 (.A0(timeout_count[27]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[28]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26433), 
          .COUT(n26434), .S0(n658[27]), .S1(n658[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_29.INIT0 = 16'h5aaa;
    defparam add_31_29.INIT1 = 16'h5aaa;
    defparam add_31_29.INJECT1_0 = "NO";
    defparam add_31_29.INJECT1_1 = "NO";
    OB Stepper_Y_M2_pad (.I(Stepper_Y_M2_c_2), .O(Stepper_Y_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    OB Stepper_Y_M1_pad (.I(Stepper_Y_M1_c_1), .O(Stepper_Y_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    CCU2D add_31_15 (.A0(timeout_count[13]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[14]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26426), 
          .COUT(n26427), .S0(n658[13]), .S1(n658[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_15.INIT0 = 16'h5aaa;
    defparam add_31_15.INIT1 = 16'h5aaa;
    defparam add_31_15.INJECT1_0 = "NO";
    defparam add_31_15.INJECT1_1 = "NO";
    OB Stepper_Y_M0_pad (.I(Stepper_Y_M0_c_0), .O(Stepper_Y_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:29])
    OB Stepper_Y_Dir_pad (.I(Stepper_Y_Dir_c), .O(Stepper_Y_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:30])
    OB Stepper_Y_Step_pad (.I(Stepper_Y_Step_c), .O(Stepper_Y_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(376[17:31])
    OB Stepper_X_En_pad (.I(Stepper_X_En_c), .O(Stepper_X_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    OB Stepper_X_M2_pad (.I(Stepper_X_M2_c_2), .O(Stepper_X_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    OB Stepper_X_M1_pad (.I(Stepper_X_M1_c_1), .O(Stepper_X_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    OB Stepper_X_M0_pad (.I(Stepper_X_M0_c_0), .O(Stepper_X_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:29])
    OB Stepper_X_Dir_pad (.I(Stepper_X_Dir_c), .O(Stepper_X_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:30])
    OB Stepper_X_Step_pad (.I(Stepper_X_Step_c), .O(Stepper_X_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(368[17:31])
    OB status_led_pad_0 (.I(VCC_net), .O(status_led[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    OB status_led_pad_1 (.I(VCC_net), .O(status_led[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    OB status_led_pad_2 (.I(VCC_net), .O(status_led[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    OB uart_tx_pad (.I(uart_tx_c), .O(uart_tx));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[14:21])
    BB expansion4_pad (.I(n11008), .T(n11007), .B(expansion4), .O(expansion4_out));
    CCU2D add_31_13 (.A0(timeout_count[11]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[12]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26425), 
          .COUT(n26426), .S0(n658[11]), .S1(n658[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_13.INIT0 = 16'h5aaa;
    defparam add_31_13.INIT1 = 16'h5aaa;
    defparam add_31_13.INJECT1_0 = "NO";
    defparam add_31_13.INJECT1_1 = "NO";
    FD1P3IX timeout_count__i1 (.D(n100_adj_1351[1]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i1.GSR = "ENABLED";
    FD1P3IX timeout_count__i2 (.D(n100_adj_1351[2]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i2.GSR = "ENABLED";
    FD1P3IX timeout_count__i3 (.D(n100_adj_1351[3]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i3.GSR = "ENABLED";
    FD1P3IX timeout_count__i4 (.D(n658[4]), .SP(n9369), .CD(n9581), .CK(debug_c_c), 
            .Q(timeout_count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i4.GSR = "ENABLED";
    FD1P3IX timeout_count__i5 (.D(n658[5]), .SP(n9369), .CD(n9581), .CK(debug_c_c), 
            .Q(timeout_count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i5.GSR = "ENABLED";
    FD1P3IX timeout_count__i6 (.D(n658[6]), .SP(n9369), .CD(n9581), .CK(debug_c_c), 
            .Q(timeout_count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i6.GSR = "ENABLED";
    FD1P3IX timeout_count__i7 (.D(n658[7]), .SP(n9369), .CD(n9581), .CK(debug_c_c), 
            .Q(timeout_count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i7.GSR = "ENABLED";
    FD1P3IX timeout_count__i8 (.D(n658[8]), .SP(n9369), .CD(n9581), .CK(debug_c_c), 
            .Q(timeout_count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i8.GSR = "ENABLED";
    FD1P3IX timeout_count__i9 (.D(n658[9]), .SP(n9369), .CD(n9581), .CK(debug_c_c), 
            .Q(timeout_count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i9.GSR = "ENABLED";
    FD1P3IX timeout_count__i10 (.D(n658[10]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i10.GSR = "ENABLED";
    FD1P3IX timeout_count__i11 (.D(n658[11]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i11.GSR = "ENABLED";
    FD1P3IX timeout_count__i12 (.D(n658[12]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i12.GSR = "ENABLED";
    FD1P3IX timeout_count__i13 (.D(n658[13]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i13.GSR = "ENABLED";
    FD1P3IX timeout_count__i14 (.D(n658[14]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i14.GSR = "ENABLED";
    FD1P3IX timeout_count__i15 (.D(n658[15]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i15.GSR = "ENABLED";
    FD1P3IX timeout_count__i16 (.D(n658[16]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i16.GSR = "ENABLED";
    FD1P3IX timeout_count__i17 (.D(n658[17]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i17.GSR = "ENABLED";
    FD1P3IX timeout_count__i18 (.D(n658[18]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i18.GSR = "ENABLED";
    FD1P3IX timeout_count__i19 (.D(n658[19]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i19.GSR = "ENABLED";
    FD1P3IX timeout_count__i20 (.D(n658[20]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i20.GSR = "ENABLED";
    FD1P3IX timeout_count__i21 (.D(n658[21]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i21.GSR = "ENABLED";
    FD1P3IX timeout_count__i22 (.D(n658[22]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i22.GSR = "ENABLED";
    FD1P3IX timeout_count__i23 (.D(n658[23]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i23.GSR = "ENABLED";
    FD1P3IX timeout_count__i24 (.D(n658[24]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i24.GSR = "ENABLED";
    FD1P3IX timeout_count__i25 (.D(n658[25]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i25.GSR = "ENABLED";
    FD1P3IX timeout_count__i26 (.D(n658[26]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i26.GSR = "ENABLED";
    FD1P3IX timeout_count__i27 (.D(n658[27]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i27.GSR = "ENABLED";
    FD1P3IX timeout_count__i28 (.D(n658[28]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i28.GSR = "ENABLED";
    FD1P3IX timeout_count__i29 (.D(n658[29]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i29.GSR = "ENABLED";
    FD1P3IX timeout_count__i30 (.D(n658[30]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i30.GSR = "ENABLED";
    FD1P3IX timeout_count__i31 (.D(n658[31]), .SP(n9369), .CD(n9581), 
            .CK(debug_c_c), .Q(timeout_count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i31.GSR = "ENABLED";
    CCU2D add_31_11 (.A0(timeout_count[9]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[10]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26424), 
          .COUT(n26425), .S0(n658[9]), .S1(n658[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_11.INIT0 = 16'h5aaa;
    defparam add_31_11.INIT1 = 16'h5aaa;
    defparam add_31_11.INJECT1_0 = "NO";
    defparam add_31_11.INJECT1_1 = "NO";
    CCU2D add_31_27 (.A0(timeout_count[25]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[26]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26432), 
          .COUT(n26433), .S0(n658[25]), .S1(n658[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_27.INIT0 = 16'h5aaa;
    defparam add_31_27.INIT1 = 16'h5aaa;
    defparam add_31_27.INJECT1_0 = "NO";
    defparam add_31_27.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_4_lut (.A(n31512), .B(register_addr[1]), .C(n31477), 
         .D(n31443), .Z(n29137)) /* synthesis lut_function=(A (B)+!A !((C (D))+!B)) */ ;
    defparam i1_2_lut_4_lut_4_lut.init = 16'h8ccc;
    LUT4 i14486_3_lut (.A(Stepper_Y_Dir_c), .B(div_factor_reg_adj_989[5]), 
         .C(register_addr[1]), .Z(n21220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i14486_3_lut.init = 16'hcaca;
    FD1P3AX reset_count_2669_2670__i2 (.D(n33692[1]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670__i2.GSR = "ENABLED";
    LUT4 i14478_3_lut (.A(Stepper_Y_En_c), .B(div_factor_reg_adj_989[6]), 
         .C(register_addr[1]), .Z(n21212)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i14478_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_281_4_lut_4_lut (.A(n31512), .B(n31477), .C(prev_select), 
         .D(n31474), .Z(n31425)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_rep_281_4_lut_4_lut.init = 16'h0400;
    LUT4 i14475_3_lut (.A(control_reg_adj_988[3]), .B(div_factor_reg_adj_989[3]), 
         .C(register_addr[1]), .Z(n21209)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i14475_3_lut.init = 16'hcaca;
    CCU2D add_31_25 (.A0(timeout_count[23]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[24]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26431), 
          .COUT(n26432), .S0(n658[23]), .S1(n658[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_25.INIT0 = 16'h5aaa;
    defparam add_31_25.INIT1 = 16'h5aaa;
    defparam add_31_25.INJECT1_0 = "NO";
    defparam add_31_25.INJECT1_1 = "NO";
    CCU2D add_31_23 (.A0(timeout_count[21]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[22]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26430), 
          .COUT(n26431), .S0(n658[21]), .S1(n658[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_23.INIT0 = 16'h5aaa;
    defparam add_31_23.INIT1 = 16'h5aaa;
    defparam add_31_23.INJECT1_0 = "NO";
    defparam add_31_23.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_511 (.A(n31512), .B(prev_select_adj_694), 
         .C(n31470), .D(select[4]), .Z(n14651)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_511.init = 16'h1000;
    FD1P3AX reset_count_2669_2670__i3 (.D(n33692[2]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670__i3.GSR = "ENABLED";
    FD1P3AX reset_count_2669_2670__i4 (.D(n33692[3]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670__i4.GSR = "ENABLED";
    FD1P3AX reset_count_2669_2670__i5 (.D(n33692[4]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670__i5.GSR = "ENABLED";
    FD1P3AX reset_count_2669_2670__i6 (.D(n33692[5]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670__i6.GSR = "ENABLED";
    FD1P3AX reset_count_2669_2670__i7 (.D(n33692[6]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670__i7.GSR = "ENABLED";
    FD1P3AX reset_count_2669_2670__i8 (.D(n33692[7]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670__i8.GSR = "ENABLED";
    FD1P3AX reset_count_2669_2670__i9 (.D(n33692[8]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670__i9.GSR = "ENABLED";
    FD1P3AX reset_count_2669_2670__i10 (.D(n33692[9]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670__i10.GSR = "ENABLED";
    FD1P3AX reset_count_2669_2670__i11 (.D(n33692[10]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670__i11.GSR = "ENABLED";
    FD1P3AX reset_count_2669_2670__i12 (.D(n33692[11]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670__i12.GSR = "ENABLED";
    FD1P3AX reset_count_2669_2670__i13 (.D(n33692[12]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670__i13.GSR = "ENABLED";
    FD1P3AX reset_count_2669_2670__i14 (.D(n33692[13]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670__i14.GSR = "ENABLED";
    FD1P3AX reset_count_2669_2670__i15 (.D(n33692[14]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670__i15.GSR = "ENABLED";
    CCU2D add_31_21 (.A0(timeout_count[19]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[20]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26429), 
          .COUT(n26430), .S0(n658[19]), .S1(n658[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_21.INIT0 = 16'h5aaa;
    defparam add_31_21.INIT1 = 16'h5aaa;
    defparam add_31_21.INJECT1_0 = "NO";
    defparam add_31_21.INJECT1_1 = "NO";
    CCU2D reset_count_2669_2670_add_4_15 (.A0(reset_count[13]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[14]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n26890), .S0(n33692[13]), .S1(n33692[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670_add_4_15.INIT0 = 16'hfaaa;
    defparam reset_count_2669_2670_add_4_15.INIT1 = 16'hfaaa;
    defparam reset_count_2669_2670_add_4_15.INJECT1_0 = "NO";
    defparam reset_count_2669_2670_add_4_15.INJECT1_1 = "NO";
    CCU2D reset_count_2669_2670_add_4_13 (.A0(reset_count[11]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[12]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n26889), .COUT(n26890), .S0(n33692[11]), .S1(n33692[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670_add_4_13.INIT0 = 16'hfaaa;
    defparam reset_count_2669_2670_add_4_13.INIT1 = 16'hfaaa;
    defparam reset_count_2669_2670_add_4_13.INJECT1_0 = "NO";
    defparam reset_count_2669_2670_add_4_13.INJECT1_1 = "NO";
    CCU2D reset_count_2669_2670_add_4_11 (.A0(reset_count[9]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[10]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n26888), .COUT(n26889), .S0(n33692[9]), .S1(n33692[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670_add_4_11.INIT0 = 16'hfaaa;
    defparam reset_count_2669_2670_add_4_11.INIT1 = 16'hfaaa;
    defparam reset_count_2669_2670_add_4_11.INJECT1_0 = "NO";
    defparam reset_count_2669_2670_add_4_11.INJECT1_1 = "NO";
    CCU2D reset_count_2669_2670_add_4_9 (.A0(reset_count[7]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[8]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n26887), .COUT(n26888), .S0(n33692[7]), .S1(n33692[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670_add_4_9.INIT0 = 16'hfaaa;
    defparam reset_count_2669_2670_add_4_9.INIT1 = 16'hfaaa;
    defparam reset_count_2669_2670_add_4_9.INJECT1_0 = "NO";
    defparam reset_count_2669_2670_add_4_9.INJECT1_1 = "NO";
    \ArmPeripheral(axis_haddr=8'b0100000)  arm_z (.read_value({read_value_adj_1030}), 
            .debug_c_c(debug_c_c), .n2847(n2847), .GND_net(battery_voltage[15]), 
            .VCC_net(VCC_net), .Stepper_Z_nFault_c(Stepper_Z_nFault_c), 
            .n31512(n31512), .\read_size[0] (read_size_adj_1031[0]), .n27753(n27753), 
            .Stepper_Z_M0_c_0(Stepper_Z_M0_c_0), .n31420(n31420), .databus({databus}), 
            .limit_latched(limit_latched_adj_702), .prev_limit_latched(prev_limit_latched_adj_703), 
            .n9305(n9305), .prev_select(prev_select_adj_738), .n31483(n31483), 
            .\read_size[2] (read_size_adj_1031[2]), .n29301(n29301), .\register_addr[1] (register_addr[1]), 
            .\register_addr[5] (register_addr[5]), .n31497(n31497), .rw(rw), 
            .\select[4] (select[4]), .n52(n52_adj_695), .\read_size[0]_adj_312 (read_size_adj_992[0]), 
            .n5(n5), .prev_select_adj_313(prev_select_adj_694), .n31422(n31422), 
            .\steps_reg[7] (steps_reg_adj_1029[7]), .n31601(n31601), .n31556(n31556), 
            .n31591(n31591), .n31596(n31596), .\register_addr[4] (register_addr[4]), 
            .n29271(n29271), .n31464(n31464), .Stepper_Z_M1_c_1(Stepper_Z_M1_c_1), 
            .\register_addr[0] (register_addr[0]), .n29235(n29235), .n31504(n31504), 
            .\read_size[2]_adj_314 (read_size_adj_980[2]), .n9(n9_adj_899), 
            .Stepper_Z_M2_c_2(Stepper_Z_M2_c_2), .n14523(n14523), .n610(n580_adj_1049[2]), 
            .n608(n580_adj_1049[4]), .Stepper_Z_Dir_c(Stepper_Z_Dir_c), 
            .Stepper_Z_En_c(Stepper_Z_En_c), .n11209(n11209), .n14547(n14547), 
            .\register_addr[3] (register_addr[3]), .\register_addr[2] (register_addr[2]), 
            .n31541(n31541), .n6(n33625[0]), .n4007(n4007), .Stepper_Z_Step_c(Stepper_Z_Step_c), 
            .limit_c_2(limit_c_2), .n11(n11), .n31411(n31411), .n16842(n16842), 
            .n8264(n8264), .n8298(n8298)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(610[25] 623[45])
    LUT4 i3_4_lut_4_lut (.A(n31512), .B(n31556), .C(n31596), .D(n29237), 
         .Z(n35)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i3_4_lut_4_lut.init = 16'h0100;
    CCU2D reset_count_2669_2670_add_4_7 (.A0(reset_count[5]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[6]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n26886), .COUT(n26887), .S0(n33692[5]), .S1(n33692[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670_add_4_7.INIT0 = 16'hfaaa;
    defparam reset_count_2669_2670_add_4_7.INIT1 = 16'hfaaa;
    defparam reset_count_2669_2670_add_4_7.INJECT1_0 = "NO";
    defparam reset_count_2669_2670_add_4_7.INJECT1_1 = "NO";
    CCU2D reset_count_2669_2670_add_4_5 (.A0(reset_count[3]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[4]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n26885), .COUT(n26886), .S0(n33692[3]), .S1(n33692[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670_add_4_5.INIT0 = 16'hfaaa;
    defparam reset_count_2669_2670_add_4_5.INIT1 = 16'hfaaa;
    defparam reset_count_2669_2670_add_4_5.INJECT1_0 = "NO";
    defparam reset_count_2669_2670_add_4_5.INJECT1_1 = "NO";
    \ArmPeripheral(axis_haddr=8'b010000)  arm_y (.debug_c_c(debug_c_c), .VCC_net(VCC_net), 
            .GND_net(battery_voltage[15]), .Stepper_Y_nFault_c(Stepper_Y_nFault_c), 
            .n31512(n31512), .n4095({n4095}), .\read_size[0] (read_size_adj_992[0]), 
            .n14651(n14651), .n27752(n27752), .Stepper_Y_M0_c_0(Stepper_Y_M0_c_0), 
            .databus({databus}), .prev_step_clk(prev_step_clk_adj_659), 
            .step_clk(step_clk_adj_658), .limit_latched(limit_latched_adj_656), 
            .prev_limit_latched(prev_limit_latched_adj_657), .n9301(n9301), 
            .prev_select(prev_select_adj_694), .n31446(n31446), .n29271(n29271), 
            .n29492(n29492), .Stepper_Y_M1_c_1(Stepper_Y_M1_c_1), .\register_addr[0] (register_addr[0]), 
            .\div_factor_reg[9] (div_factor_reg_adj_989[9]), .\div_factor_reg[6] (div_factor_reg_adj_989[6]), 
            .\div_factor_reg[5] (div_factor_reg_adj_989[5]), .\div_factor_reg[4] (div_factor_reg_adj_989[4]), 
            .\div_factor_reg[3] (div_factor_reg_adj_989[3]), .\control_reg[7] (control_reg_adj_988[7]), 
            .n12149(n12149), .Stepper_Y_En_c(Stepper_Y_En_c), .Stepper_Y_Dir_c(Stepper_Y_Dir_c), 
            .\control_reg[4] (control_reg_adj_988[4]), .\control_reg[3] (control_reg_adj_988[3]), 
            .Stepper_Y_M2_c_2(Stepper_Y_M2_c_2), .\read_size[2] (read_size_adj_992[2]), 
            .n29200(n29200), .\steps_reg[9] (steps_reg_adj_990[9]), .\steps_reg[6] (steps_reg_adj_990[6]), 
            .\steps_reg[5] (steps_reg_adj_990[5]), .\steps_reg[4] (steps_reg_adj_990[4]), 
            .\steps_reg[3] (steps_reg_adj_990[3]), .read_value({read_value_adj_991}), 
            .n9548(n9548), .\register_addr[1] (register_addr[1]), .n29113(n29113), 
            .limit_c_1(limit_c_1), .int_step(int_step), .n22(n22), .n31419(n31419), 
            .n29114(n29114), .n21214(n21214), .n21222(n21222), .n28827(n28827), 
            .n6808(n6779[3]), .n32(n32_adj_619), .n27484(n27484), .n224({n224_adj_995}), 
            .n8636(n8635[7]), .n8194(n8194), .n31408(n31408), .n16841(n16841), 
            .n8160(n8160)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(595[25] 608[45])
    CCU2D reset_count_2669_2670_add_4_3 (.A0(reset_count[1]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[2]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n26884), .COUT(n26885), .S0(n33692[1]), .S1(n33692[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670_add_4_3.INIT0 = 16'hfaaa;
    defparam reset_count_2669_2670_add_4_3.INIT1 = 16'hfaaa;
    defparam reset_count_2669_2670_add_4_3.INJECT1_0 = "NO";
    defparam reset_count_2669_2670_add_4_3.INJECT1_1 = "NO";
    CCU2D reset_count_2669_2670_add_4_1 (.A0(battery_voltage[15]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[0]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .COUT(n26884), .S1(n33692[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2669_2670_add_4_1.INIT0 = 16'hF000;
    defparam reset_count_2669_2670_add_4_1.INIT1 = 16'h0555;
    defparam reset_count_2669_2670_add_4_1.INJECT1_0 = "NO";
    defparam reset_count_2669_2670_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(register_addr[1]), .B(n9548), .Z(n29113)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_2_lut.init = 16'h2222;
    RCPeripheral rc_receiver (.n2(n2_adj_925), .databus({databus}), .\read_value[10] (read_value_adj_1069[10]), 
            .n8(n8_adj_927), .n31426(n31426), .\register_addr[0] (register_addr[0]), 
            .read_value({read_value}), .read_value_adj_308({read_value_adj_979}), 
            .n46(n46), .n52(n52), .databus_out({databus_out}), .rw(rw), 
            .read_value_adj_309({read_value_adj_991}), .\read_value[10]_adj_157 (read_value_adj_1115[10]), 
            .n52_adj_158(n52_adj_695), .n31447(n31447), .n2_adj_159(n2_adj_929), 
            .\read_value[9]_adj_160 (read_value_adj_1069[9]), .n8_adj_161(n8_adj_931), 
            .\read_value[9]_adj_162 (read_value_adj_1115[9]), .n2_adj_163(n2_adj_926), 
            .\select[7] (select[7]), .n176(n176), .\read_value[8]_adj_164 (read_value_adj_1069[8]), 
            .n8_adj_165(n8_adj_928), .\register_addr[1] (register_addr[1]), 
            .n2_adj_166(n2_adj_937), .\read_value[24]_adj_167 (read_value_adj_1069[24]), 
            .n8_adj_168(n8), .\read_value[24]_adj_169 (read_value_adj_1115[24]), 
            .\read_value[8]_adj_170 (read_value_adj_1115[8]), .n2_adj_171(n2_adj_930), 
            .\read_value[7]_adj_172 (read_value_adj_1115[7]), .\read_value[7]_adj_173 (read_value_adj_1107[7]), 
            .n31444(n31444), .n3(n3_adj_932), .read_value_adj_310({read_value_adj_972}), 
            .n64(n64), .n66(n66), .read_value_adj_311({read_value_adj_1131}), 
            .\read_value[14]_adj_190 (read_value_adj_1115[14]), .n2_adj_191(n2_adj_741), 
            .\read_value[6]_adj_192 (read_value_adj_1115[6]), .\read_value[6]_adj_193 (read_value_adj_1107[6]), 
            .n3_adj_194(n3_adj_948), .n2_adj_195(n2_adj_606), .\read_value[5]_adj_196 (read_value_adj_1115[5]), 
            .\read_value[5]_adj_197 (read_value_adj_1107[5]), .n33385(n33385), 
            .n3_adj_198(n3), .n2_adj_199(n2_adj_902), .\read_value[4]_adj_200 (read_value_adj_1115[4]), 
            .\read_value[4]_adj_201 (read_value_adj_1107[4]), .n3_adj_202(n3_adj_901), 
            .n2_adj_203(n2_adj_817), .\read_value[3]_adj_204 (read_value_adj_1115[3]), 
            .\read_value[3]_adj_205 (read_value_adj_1107[3]), .n2_adj_206(n2_adj_900), 
            .\read_value[22]_adj_207 (read_value_adj_1069[22]), .n8_adj_208(n8_adj_740), 
            .n3_adj_209(n3_adj_947), .n2_adj_210(n2_adj_936), .\read_value[2]_adj_211 (read_value_adj_1115[2]), 
            .\read_value[2]_adj_212 (read_value_adj_1107[2]), .\read_value[22]_adj_213 (read_value_adj_1115[22]), 
            .n3_adj_214(n3_adj_620), .n10(n10), .\read_value[1]_adj_215 (read_value_adj_1107[1]), 
            .n3_adj_216(n3_adj_701), .\read_value[1]_adj_217 (read_value_adj_1069[1]), 
            .n2_adj_218(n2_adj_923), .\read_value[13]_adj_219 (read_value_adj_1069[13]), 
            .n8_adj_220(n8_adj_924), .n2_adj_221(n2_adj_742), .\read_value[13]_adj_222 (read_value_adj_1115[13]), 
            .\read_value[23]_adj_223 (read_value_adj_1069[23]), .n8_adj_224(n8_adj_739), 
            .n2_adj_225(n2_adj_700), .n2_adj_226(n2_adj_933), .\read_value[12]_adj_227 (read_value_adj_1069[12]), 
            .n8_adj_228(n8_adj_935), .\read_value[23]_adj_229 (read_value_adj_1115[23]), 
            .\read_value[12]_adj_230 (read_value_adj_1115[12]), .\read_value[21]_adj_231 (read_value_adj_1069[21]), 
            .n8_adj_232(n8_adj_945), .read_size({read_size}), .\select[1] (select[1]), 
            .n13(n13_adj_699), .n31483(n31483), .n9(n9), .\read_size[0]_adj_233 (read_size_adj_1031[0]), 
            .n18(n18), .\read_size[0]_adj_234 (read_size_adj_1108[0]), .\read_size[0]_adj_235 (read_size_adj_973[0]), 
            .n31465(n31465), .\select[2] (select[2]), .n14(n14_adj_698), 
            .n31474(n31474), .n5(n5), .\read_size[0]_adj_236 (read_size_adj_980[0]), 
            .\read_size[0]_adj_237 (read_size_adj_1132[0]), .n31445(n31445), 
            .\select[5] (select[5]), .\read_size[0]_adj_238 (read_size_adj_1070[0]), 
            .n2_adj_239(n2), .\read_value[11]_adj_240 (read_value_adj_1069[11]), 
            .n8_adj_241(n8_adj_608), .n6(n6), .\read_size[2]_adj_242 (read_size_adj_1070[2]), 
            .\reg_size[2] (reg_size[2]), .\read_size[2]_adj_243 (read_size_adj_1031[2]), 
            .n9_adj_244(n9_adj_899), .\read_size[2]_adj_245 (read_size_adj_1116[2]), 
            .n31471(n31471), .\read_value[11]_adj_246 (read_value_adj_1115[11]), 
            .\read_value[21]_adj_247 (read_value_adj_1115[21]), .n2_adj_248(n2_adj_609), 
            .\read_value[25]_adj_249 (read_value_adj_1069[25]), .n8_adj_250(n8_adj_697), 
            .\read_value[25]_adj_251 (read_value_adj_1115[25]), .\register_addr[2] (register_addr[2]), 
            .n2_adj_252(n2_adj_942), .n2_adj_253(n2_adj_915), .\read_value[20]_adj_254 (read_value_adj_1069[20]), 
            .n8_adj_255(n8_adj_946), .\read_value[16]_adj_256 (read_value_adj_1069[16]), 
            .n8_adj_257(n8_adj_916), .n31588(n31588), .\sendcount[1] (sendcount[1]), 
            .n13156(n13156), .n31457(n31457), .\read_value[20]_adj_258 (read_value_adj_1115[20]), 
            .n2_adj_259(n2_adj_921), .n2_adj_260(n2_adj_605), .\read_value[0]_adj_261 (read_value_adj_1115[0]), 
            .\read_value[0]_adj_262 (read_value_adj_1107[0]), .n3_adj_263(n3_adj_607), 
            .n2_adj_264(n2_adj_914), .\read_value[26]_adj_265 (read_value_adj_1069[26]), 
            .n8_adj_266(n8_adj_913), .\read_value[26]_adj_267 (read_value_adj_1115[26]), 
            .\read_value[16]_adj_268 (read_value_adj_1115[16]), .n2_adj_269(n2_adj_943), 
            .\read_value[19]_adj_270 (read_value_adj_1069[19]), .n8_adj_271(n8_adj_818), 
            .n29237(n29237), .n2_adj_272(n2_adj_918), .\read_value[19]_adj_273 (read_value_adj_1115[19]), 
            .n2_adj_274(n2_adj_934), .\read_value[18]_adj_275 (read_value_adj_1069[18]), 
            .n8_adj_276(n8_adj_813), .n2_adj_277(n2_adj_903), .\read_value[31]_adj_278 (read_value_adj_1069[31]), 
            .n8_adj_279(n8_adj_904), .\read_value[14]_adj_280 (read_value_adj_1069[14]), 
            .n8_adj_281(n8_adj_922), .\read_value[31]_adj_282 (read_value_adj_1115[31]), 
            .n2_adj_283(n2_adj_816), .\read_value[30]_adj_284 (read_value_adj_1069[30]), 
            .n8_adj_285(n8_adj_906), .\read_value[18]_adj_286 (read_value_adj_1115[18]), 
            .\read_value[30]_adj_287 (read_value_adj_1115[30]), .n2_adj_288(n2_adj_908), 
            .\read_value[17]_adj_289 (read_value_adj_1115[17]), .\read_value[29]_adj_290 (read_value_adj_1069[29]), 
            .n8_adj_291(n8_adj_815), .\read_value[29]_adj_292 (read_value_adj_1115[29]), 
            .n2_adj_293(n2_adj_911), .n2_adj_294(n2_adj_917), .\read_value[15]_adj_295 (read_value_adj_1069[15]), 
            .n8_adj_296(n8_adj_920), .\read_value[28]_adj_297 (read_value_adj_1069[28]), 
            .n8_adj_298(n8_adj_909), .\read_value[17]_adj_299 (read_value_adj_1069[17]), 
            .n8_adj_300(n8_adj_919), .\read_value[28]_adj_301 (read_value_adj_1115[28]), 
            .n2_adj_302(n2_adj_912), .\read_value[27]_adj_303 (read_value_adj_1069[27]), 
            .n8_adj_304(n8_adj_814), .\read_value[15]_adj_305 (read_value_adj_1115[15]), 
            .\read_value[27]_adj_306 (read_value_adj_1115[27]), .GND_net(battery_voltage[15]), 
            .debug_c_c(debug_c_c), .n33387(n33387), .rc_ch8_c(rc_ch8_c), 
            .n29818(n29818), .n33386(n33386), .n13957(n13957), .n27564(n27564), 
            .n29784(n29784), .rc_ch7_c(rc_ch7_c), .n33388(n33388), .n27543(n27543), 
            .n29827(n29827), .rc_ch4_c(rc_ch4_c), .n27550(n27550), .n29838(n29838), 
            .rc_ch3_c(rc_ch3_c), .n14500(n14500), .n27541(n27541), .n29840(n29840), 
            .n29530(n29530), .n29944(n29944), .n14_adj_307(n14_adj_910), 
            .n29832(n29832), .rc_ch2_c(rc_ch2_c), .n31412(n31412), .n14513(n14513), 
            .n29847(n29847), .n27536(n27536), .n31512(n31512), .n14514(n14514), 
            .rc_ch1_c(rc_ch1_c), .n29830(n29830), .n27547(n27547), .n29811(n29811)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(708[15] 720[41])
    LUT4 i15746_1_lut_rep_471 (.A(reset_count[14]), .B(reset_count[12]), 
         .C(reset_count[13]), .D(n29264), .Z(n33390)) /* synthesis lut_function=(!(A+(B (C)+!B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam i15746_1_lut_rep_471.init = 16'h0515;
    SabertoothSerialPeripheral motor_serial (.\read_size[0] (read_size_adj_973[0]), 
            .debug_c_c(debug_c_c), .n9379(n9379), .n13908(n13908), .n31512(n31512), 
            .\databus[0] (databus[0]), .\select[2] (select[2]), .read_value({read_value_adj_972}), 
            .n9542(n9542), .rw(rw), .n64(n64), .n31601(n31601), .\register[0][7] (\register[0]_adj_971 [7]), 
            .n31582(n31582), .\reset_count[14] (reset_count[14]), .n22484(n22484), 
            .n11236(n11236), .\databus[7] (databus[7]), .\databus[6] (databus[6]), 
            .\databus[5] (databus[5]), .\databus[4] (databus[4]), .\databus[3] (databus[3]), 
            .\databus[2] (databus[2]), .\databus[1] (databus[1]), .\register_addr[0] (register_addr[0]), 
            .n31413(n31413), .GND_net(battery_voltage[15]), .n1156(n1156), 
            .n31537(n31537), .\reset_count[8] (reset_count[8]), .\reset_count[7] (reset_count[7]), 
            .n29332(n29332), .state({state_adj_1308}), .n29170(n29170), 
            .n31596(n31596), .n31556(n31556), .n31576(n31576), .n9(n9_adj_938), 
            .n33385(n33385), .n31443(n31443), .n31590(n31590), .n35(n35), 
            .n4181(n4181), .\register_addr[5] (register_addr[5]), .n31464(n31464), 
            .n13917(n13917), .\reset_count[11] (reset_count[11]), .n21503(n21503), 
            .n27250(n27250), .n29264(n29264), .n14783(n14783), .n31530(n31530), 
            .n9297(n9297), .n31463(n31463), .n11073(n11073), .n8507(n8507), 
            .n29786(n29786), .select_clk(select_clk), .n2967(n2967), .n107(n107)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(530[29] 538[56])
    GSR GSR_INST (.GSR(VCC_net));
    LUT4 Select_4241_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[24]), 
         .D(rw), .Z(n8)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4241_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    \ProtocolInterface(baud_div=12)  protocol_interface (.register_addr({Open_0, 
            Open_1, register_addr[5:0]}), .debug_c_c(debug_c_c), .databus({databus}), 
            .\select[7] (select[7]), .n33390(n33390), .\select[5] (select[5]), 
            .\select[4] (select[4]), .\select[3] (select[3]), .\select[2] (select[2]), 
            .\select[1] (select[1]), .databus_out({databus_out}), .n13834(n13834), 
            .\sendcount[1] (sendcount[1]), .n31556(n31556), .n29301(n29301), 
            .n31533(n31533), .n29200(n29200), .debug_c_5(debug_c_5), .n31497(n31497), 
            .rw(rw), .n31426(n31426), .prev_select(prev_select_adj_780), 
            .n31428(n31428), .n31596(n31596), .n31470(n31470), .n31466(n31466), 
            .n31427(n31427), .\register[1][19] (\register[1]_adj_1105 [19]), 
            .n59(n99_adj_1332[19]), .n31501(n31501), .\register[1][20] (\register[1]_adj_1105 [20]), 
            .n57(n99_adj_1332[20]), .\register[1][26] (\register[1]_adj_1105 [26]), 
            .n45(n99_adj_1332[26]), .force_pause(force_pause), .\register[2] ({\register[2] }), 
            .\register[1][0] (\register[1]_adj_1105 [0]), .n97(n99_adj_1332[0]), 
            .n31504(n31504), .prev_select_adj_5(prev_select), .n31512(n31512), 
            .n13941(n13941), .n1492(n1474[14]), .n29170(n29170), .n29295(n29295), 
            .n29069(n29069), .n29293(n29293), .n31436(n31436), .n303(n303), 
            .n56(n56), .n29294(n29294), .n29066(n29066), .n29056(n29056), 
            .n29053(n29053), .n29065(n29065), .n29063(n29063), .n29050(n29050), 
            .n224({n224_adj_1073}), .n3922({n3922}), .n29052(n29052), 
            .n29054(n29054), .n27752(n27752), .n29067(n29067), .n29057(n29057), 
            .n29068(n29068), .n29071(n29071), .n29072(n29072), .n27753(n27753), 
            .n29070(n29070), .n29058(n29058), .n29059(n29059), .n29064(n29064), 
            .n29060(n29060), .n29258(n29258), .n29062(n29062), .n29055(n29055), 
            .n29051(n29051), .n29049(n29049), .n29061(n29061), .n29048(n29048), 
            .prev_select_adj_6(prev_select_adj_738), .n2847(n2847), .n66(n66), 
            .\register[0][2] (\register[0] [2]), .read_value({read_value_adj_1030}), 
            .n33385(n33385), .n2(n2_adj_742), .n31465(n31465), .n2_adj_7(n2_adj_900), 
            .n2_adj_8(n2_adj_700), .n2_adj_9(n2_adj_942), .n2_adj_10(n2_adj_609), 
            .n31541(n31541), .n31450(n31450), .n31478(n31478), .n31471(n31471), 
            .n2_adj_11(n2_adj_937), .n2_adj_12(n2_adj_943), .n2_adj_13(n2_adj_934), 
            .n31474(n31474), .n2_adj_14(n2_adj_917), .n2_adj_15(n2_adj_915), 
            .n2_adj_16(n2_adj_918), .n2_adj_17(n2_adj_921), .n2_adj_18(n2_adj_923), 
            .n2_adj_19(n2_adj_933), .n2_adj_20(n2), .n2_adj_21(n2_adj_925), 
            .n2_adj_22(n2_adj_929), .n2_adj_23(n2_adj_926), .n3(n3_adj_932), 
            .n3_adj_24(n3_adj_948), .n3_adj_25(n3), .n31590(n31590), .n31477(n31477), 
            .n3_adj_26(n3_adj_901), .n3_adj_27(n3_adj_947), .n3_adj_28(n3_adj_620), 
            .n3_adj_29(n3_adj_701), .n3_adj_30(n3_adj_607), .n2_adj_31(n2_adj_903), 
            .n2_adj_32(n2_adj_816), .n2_adj_33(n2_adj_908), .n2_adj_34(n2_adj_911), 
            .n2_adj_35(n2_adj_912), .n2_adj_36(n2_adj_914), .n31483(n31483), 
            .n14454(n14454), .n9538(n9538), .n35(n35), .n27465(n27465), 
            .n33384(n33384), .n31446(n31446), .debug_c_7(debug_c_7), .\read_size[2] (read_size_adj_992[2]), 
            .n29235(n29235), .n31445(n31445), .n52(n52), .n31443(n31443), 
            .n29237(n29237), .n176(n176), .n31449(n31449), .n31571(n31571), 
            .n16013(n16013), .n31457(n31457), .n31582(n31582), .n13908(n13908), 
            .n11236(n11236), .n31435(n31435), .n30306(n30306), .n29221(n29221), 
            .n31526(n31526), .n31420(n31420), .n30304(n30304), .\control_reg[7] (control_reg[7]), 
            .n1(n1), .n31530(n31530), .n31540(n31540), .n13156(n13156), 
            .n13(n13_adj_699), .n18(n18), .n14(n14_adj_698), .\reg_size[2] (reg_size[2]), 
            .n31588(n31588), .n31591(n31591), .n27442(n27442), .\control_reg[7]_adj_37 (control_reg_adj_1066[7]), 
            .n31601(n31601), .n32(n32), .n4(n4), .n5834(n5834), .prev_select_adj_38(prev_select_adj_898), 
            .\reset_count[14] (reset_count[14]), .n22484(n22484), .n2870(n2870), 
            .n224_adj_91({n224_adj_995}), .n4095({n4095}), .n31576(n31576), 
            .\read_value[7]_adj_71 (read_value_adj_1069[7]), .n2_adj_72(n2_adj_930), 
            .\read_value[5]_adj_73 (read_value_adj_1069[5]), .n2_adj_74(n2_adj_606), 
            .n31473(n31473), .\read_value[4]_adj_75 (read_value_adj_1069[4]), 
            .n2_adj_76(n2_adj_902), .\read_value[6]_adj_77 (read_value_adj_1069[6]), 
            .n2_adj_78(n2_adj_741), .\read_value[3]_adj_79 (read_value_adj_1069[3]), 
            .n2_adj_80(n2_adj_817), .\read_value[2]_adj_81 (read_value_adj_1069[2]), 
            .n2_adj_82(n2_adj_936), .\read_value[0]_adj_83 (read_value_adj_1069[0]), 
            .n2_adj_84(n2_adj_605), .n27445(n27445), .n34(n34), .n29257(n29257), 
            .n9331(n9331), .n1486(n1474[20]), .\register[0][5] (\register[0]_adj_1130 [5]), 
            .expansion5_c(expansion5_c), .\register[1][5] (\register[1]_adj_1129 [5]), 
            .debug_c_2(debug_c_2), .n1489(n1474[17]), .debug_c_3(debug_c_3), 
            .n9379(n9379), .n29492(n29492), .prev_select_adj_85(prev_select_adj_694), 
            .\steps_reg[7] (steps_reg_adj_1029[7]), .n11(n11), .debug_c_4(debug_c_4), 
            .n31502(n31502), .n6006(n5974[0]), .\steps_reg[5] (steps_reg_adj_990[5]), 
            .n14_adj_86(n14), .\register[0][4] (\register[0]_adj_1130 [4]), 
            .expansion4_out(expansion4_out), .\register[1][4] (\register[1]_adj_1129 [4]), 
            .timeout_pause(timeout_pause), .\steps_reg[6] (steps_reg_adj_990[6]), 
            .n13_adj_87(n13), .\register[0][7] (\register[0]_adj_971 [7]), 
            .n31537(n31537), .clk_1Hz(clk_1Hz), .signal_light_c(signal_light_c), 
            .\steps_reg[3] (steps_reg_adj_990[3]), .n12(n12), .\control_reg[4] (control_reg_adj_988[4]), 
            .\div_factor_reg[4] (div_factor_reg_adj_989[4]), .\steps_reg[4] (steps_reg_adj_990[4]), 
            .\control_reg[7]_adj_88 (control_reg_adj_988[7]), .n8636(n8635[7]), 
            .n13948(n13948), .n12369(n12369), .n9301(n9301), .n14523(n14523), 
            .n4007(n4007), .n31407(n31407), .n27680(n27680), .n27484(n27484), 
            .n32_adj_89(n32_adj_619), .n16765(n16765), .n9(n9_adj_938), 
            .n9305(n9305), .prev_select_adj_90(prev_select_adj_853), .n16764(n16764), 
            .n6003(n5974[3]), .n27428(n27428), .n28827(n28827), .n8654(n8653[7]), 
            .\state[3] (state_adj_1308[3]), .\state[1] (state_adj_1308[1]), 
            .\state[0] (state_adj_1308[0]), .n1156(n1156), .n73(n73), 
            .\reset_count[7] (reset_count[7]), .\reset_count[6] (reset_count[6]), 
            .\reset_count[5] (reset_count[5]), .n27250(n27250), .uart_tx_c(uart_tx_c), 
            .GND_net(battery_voltage[15]), .uart_rx_c(uart_rx_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(493[26] 503[57])
    CCU2D add_31_19 (.A0(timeout_count[17]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[18]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n26428), 
          .COUT(n26429), .S0(n658[17]), .S1(n658[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_19.INIT0 = 16'h5aaa;
    defparam add_31_19.INIT1 = 16'h5aaa;
    defparam add_31_19.INJECT1_0 = "NO";
    defparam add_31_19.INJECT1_1 = "NO";
    LUT4 Select_4238_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[25]), 
         .D(rw), .Z(n8_adj_697)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4238_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4244_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[23]), 
         .D(rw), .Z(n8_adj_739)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4244_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4247_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[22]), 
         .D(rw), .Z(n8_adj_740)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4247_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4250_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[21]), 
         .D(rw), .Z(n8_adj_945)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4250_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2658_1_lut (.A(n7847), .Z(n9369)) /* synthesis lut_function=(!(A)) */ ;
    defparam i2658_1_lut.init = 16'h5555;
    LUT4 i30_2_lut (.A(uart_rx_c), .B(prev_uart_rx), .Z(n9581)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(475[7:30])
    defparam i30_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_512 (.A(div_factor_reg_adj_989[9]), .B(n29113), .C(steps_reg_adj_990[9]), 
         .D(register_addr[0]), .Z(n29114)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_4_lut_adj_512.init = 16'hc088;
    LUT4 Select_4253_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[20]), 
         .D(rw), .Z(n8_adj_946)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4253_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4256_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[19]), 
         .D(rw), .Z(n8_adj_818)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4256_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    PFUMX i14488 (.BLUT(n21220), .ALUT(n14), .C0(register_addr[0]), .Z(n21222));
    LUT4 Select_4259_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[18]), 
         .D(rw), .Z(n8_adj_813)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4259_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4262_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[17]), 
         .D(rw), .Z(n8_adj_919)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4262_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4265_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[16]), 
         .D(rw), .Z(n8_adj_916)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4265_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i22315_2_lut (.A(int_step), .B(control_reg_adj_988[3]), .Z(Stepper_Y_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i22315_2_lut.init = 16'h9999;
    LUT4 Select_4268_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[15]), 
         .D(rw), .Z(n8_adj_920)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4268_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    PFUMX i14480 (.BLUT(n21212), .ALUT(n13), .C0(register_addr[0]), .Z(n21214));
    LUT4 Select_4271_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[14]), 
         .D(n33385), .Z(n8_adj_922)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4271_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    GlobalControlPeripheral global_control (.\register[2] ({\register[2] }), 
            .GND_net(battery_voltage[15]), .force_pause(force_pause), .debug_c_c(debug_c_c), 
            .n31512(n31512), .\databus[1] (databus[1]), .n9484(n9484), 
            .read_size({read_size}), .n14454(n14454), .n31450(n31450), 
            .prev_clk_1Hz(prev_clk_1Hz), .clk_1Hz(clk_1Hz), .\register[0][2] (\register[0] [2]), 
            .\select[1] (select[1]), .read_value({read_value}), .n29069(n29069), 
            .rw(rw), .n46(n46), .n29293(n29293), .n31478(n31478), .n29294(n29294), 
            .n29295(n29295), .n30306(n30306), .n30304(n30304), .\reset_count[14] (reset_count[14]), 
            .n22484(n22484), .xbee_pause_c(xbee_pause_c), .\register_addr[1] (register_addr[1]), 
            .\register_addr[0] (register_addr[0]), .n29170(n29170), .n9538(n9538), 
            .n6003(n5974[3]), .n29066(n29066), .n29056(n29056), .n29053(n29053), 
            .n16765(n16765), .n27428(n27428), .n29065(n29065), .n16764(n16764), 
            .n29063(n29063), .n29050(n29050), .n29052(n29052), .n29054(n29054), 
            .n29067(n29067), .n29057(n29057), .n29068(n29068), .n29071(n29071), 
            .n29072(n29072), .n29070(n29070), .n6006(n5974[0]), .n29058(n29058), 
            .n29059(n29059), .n29064(n29064), .n29060(n29060), .n29062(n29062), 
            .n29055(n29055), .n29051(n29051), .n29049(n29049), .n29061(n29061), 
            .n29048(n29048), .n29789(n29789), .n2876(n2876)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(514[45] 525[74])
    ClockDivider_U10 pwm_clk_div (.clk_255kHz(clk_255kHz), .debug_c_c(debug_c_c), 
            .n241(n241), .GND_net(battery_voltage[15]), .n7917(n7917), 
            .n31512(n31512), .n7882(n7882), .n29832(n29832), .n14513(n14513), 
            .n29830(n29830), .n14514(n14514), .n2824(n2824), .n29840(n29840), 
            .n27541(n27541), .n29847(n29847), .n27536(n27536), .n29818(n29818), 
            .n13957(n13957), .n29530(n29530), .n14(n14_adj_910), .n29944(n29944), 
            .n14500(n14500), .n29784(n29784), .n27564(n27564), .n29811(n29811), 
            .n27547(n27547), .n29827(n29827), .n27543(n27543), .n29838(n29838), 
            .n27550(n27550)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(540[15] 543[41])
    LUT4 Select_4274_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[13]), 
         .D(rw), .Z(n8_adj_924)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4274_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    PFUMX i14477 (.BLUT(n21209), .ALUT(n12), .C0(register_addr[0]), .Z(n6779[3]));
    LUT4 Select_4277_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[12]), 
         .D(rw), .Z(n8_adj_935)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4277_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4280_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[11]), 
         .D(rw), .Z(n8_adj_608)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4280_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    \ArmPeripheral(axis_haddr=8'b0)  arm_x (.debug_c_c(debug_c_c), .n31512(n31512), 
            .databus({databus}), .n4181(n4181), .\read_size[0] (read_size_adj_980[0]), 
            .n13941(n13941), .n9379(n9379), .Stepper_X_M0_c_0(Stepper_X_M0_c_0), 
            .n13917(n13917), .prev_step_clk(prev_step_clk), .step_clk(step_clk), 
            .limit_latched(limit_latched), .prev_limit_latched(prev_limit_latched), 
            .n9297(n9297), .prev_select(prev_select), .n31474(n31474), 
            .\register_addr[1] (register_addr[1]), .Stepper_X_Dir_c(Stepper_X_Dir_c), 
            .\register_addr[0] (register_addr[0]), .n1(n1), .Stepper_X_En_c(Stepper_X_En_c), 
            .Stepper_X_M1_c_1(Stepper_X_M1_c_1), .\control_reg[7] (control_reg[7]), 
            .n12159(n12159), .Stepper_X_M2_c_2(Stepper_X_M2_c_2), .\read_size[2] (read_size_adj_980[2]), 
            .n31435(n31435), .n34(n34), .n27445(n27445), .n29137(n29137), 
            .limit_c_0(limit_c_0), .read_value({read_value_adj_979}), .n31425(n31425), 
            .n24(n24), .n31421(n31421), .VCC_net(VCC_net), .GND_net(battery_voltage[15]), 
            .Stepper_X_nFault_c(Stepper_X_nFault_c), .Stepper_X_Step_c(Stepper_X_Step_c), 
            .n31409(n31409), .n8056(n8056), .n8090(n8090), .n17035(n17035)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(580[25] 593[45])
    LUT4 Select_4283_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[10]), 
         .D(n33385), .Z(n8_adj_927)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4283_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_4_lut (.A(n31512), .B(n303), .C(n31449), .D(n31571), 
         .Z(n24146)) /* synthesis lut_function=(!(A+!(B (D)+!B (C (D))))) */ ;
    defparam i2_4_lut_4_lut.init = 16'h5400;
    LUT4 Select_4286_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[9]), 
         .D(n33385), .Z(n8_adj_931)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4286_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_4_lut_adj_513 (.A(n31512), .B(n31533), .C(n31540), .D(n31422), 
         .Z(n9548)) /* synthesis lut_function=(!(A+!(B (D)+!B !(C+!(D))))) */ ;
    defparam i2_4_lut_4_lut_adj_513.init = 16'h4500;
    LUT4 Select_4289_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[8]), 
         .D(n33385), .Z(n8_adj_928)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4289_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4220_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[31]), 
         .D(n33385), .Z(n8_adj_904)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4220_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    EncoderPeripheral right_encoder (.\register_addr[0] (register_addr[0]), 
            .n31432(n31432), .prev_select(prev_select_adj_888), .debug_c_c(debug_c_c), 
            .n31471(n31471), .\read_size[0] (read_size_adj_1116[0]), .n15087(n15087), 
            .n6(n33625[0]), .encoder_rb_c(encoder_rb_c), .encoder_ra_c(encoder_ra_c), 
            .read_value({read_value_adj_1115}), .\read_size[2] (read_size_adj_1116[2]), 
            .n31541(n31541), .encoder_ri_c(encoder_ri_c), .qreset(qreset), 
            .VCC_net(VCC_net), .GND_net(battery_voltage[15]), .\quadA_delayed[1] (quadA_delayed_adj_1219[1]), 
            .n13939(n13939), .n6_adj_4(n6_adj_944), .\quadB_delayed[1] (quadB_delayed_adj_1220[1])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(682[20] 692[47])
    \ClockDividerP_SP(factor=120000)  clk_100Hz_divider (.n29792(n29792), 
            .debug_c_0(debug_c_0), .debug_c_c(debug_c_c), .n31512(n31512), 
            .n2861(n2861), .GND_net(battery_voltage[15])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(643[29] 645[61])
    LUT4 Select_4223_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[30]), 
         .D(n33385), .Z(n8_adj_906)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4223_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 m1_lut (.Z(n33384)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    LUT4 i15736_4_lut (.A(n22390), .B(n13316), .C(n21503), .D(n29332), 
         .Z(n22484)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i15736_4_lut.init = 16'hfcec;
    LUT4 i15647_3_lut (.A(reset_count[5]), .B(reset_count[6]), .C(reset_count[4]), 
         .Z(n22390)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i15647_3_lut.init = 16'hc8c8;
    LUT4 Select_4226_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[29]), 
         .D(n33385), .Z(n8_adj_815)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4226_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    EncoderPeripheral_U11 left_encoder (.\read_size[0] (read_size_adj_1108[0]), 
            .debug_c_c(debug_c_c), .n14146(n14146), .n31427(n31427), .n31450(n31450), 
            .prev_select(prev_select_adj_853), .n31465(n31465), .\read_size[2] (read_size_adj_1108[2]), 
            .n31478(n31478), .read_value({read_value_adj_1107}), .\register_addr[0] (register_addr[0]), 
            .encoder_la_c(encoder_la_c), .encoder_lb_c(encoder_lb_c), .n59(n99_adj_1332[19]), 
            .n57(n99_adj_1332[20]), .n45(n99_adj_1332[26]), .\quadA_delayed[1] (quadA_delayed_adj_1219[1]), 
            .qreset(qreset), .n6(n6_adj_944), .\quadB_delayed[1] (quadB_delayed_adj_1220[1]), 
            .n13939(n13939), .n97(n99_adj_1332[0]), .encoder_li_c(encoder_li_c), 
            .GND_net(battery_voltage[15]), .\register[1][0] (\register[1]_adj_1105 [0]), 
            .VCC_net(VCC_net), .\register[1][19] (\register[1]_adj_1105 [19]), 
            .\register[1][20] (\register[1]_adj_1105 [20]), .\register[1][26] (\register[1]_adj_1105 [26])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(671[20] 681[47])
    \ArmPeripheral(axis_haddr=8'b0110000)  arm_a (.read_value({read_value_adj_1069}), 
            .debug_c_c(debug_c_c), .n2858(n2858), .n31512(n31512), .n3922({n3922}), 
            .VCC_net(VCC_net), .GND_net(battery_voltage[15]), .Stepper_A_nFault_c(Stepper_A_nFault_c), 
            .\read_size[0] (read_size_adj_1070[0]), .n29258(n29258), .Stepper_A_M0_c_0(Stepper_A_M0_c_0), 
            .databus({databus}), .limit_latched(limit_latched_adj_744), 
            .prev_limit_latched(prev_limit_latched_adj_745), .n9331(n9331), 
            .prev_select(prev_select_adj_780), .n31445(n31445), .Stepper_A_M1_c_1(Stepper_A_M1_c_1), 
            .\register_addr[0] (register_addr[0]), .\register_addr[1] (register_addr[1]), 
            .n224({n224_adj_1073}), .n32(n32), .n32_adj_1(n32_adj_619), 
            .prev_step_clk(prev_step_clk_adj_659), .step_clk(step_clk_adj_658), 
            .n31419(n31419), .n22(n22), .prev_step_clk_adj_2(prev_step_clk), 
            .n34(n34), .step_clk_adj_3(step_clk), .n31421(n31421), .n24(n24), 
            .n31428(n31428), .\register_addr[5] (register_addr[5]), .n31497(n31497), 
            .n29271(n29271), .n31576(n31576), .n27442(n27442), .\read_size[2] (read_size_adj_1070[2]), 
            .n29257(n29257), .Stepper_A_M2_c_2(Stepper_A_M2_c_2), .Stepper_A_Dir_c(Stepper_A_Dir_c), 
            .Stepper_A_En_c(Stepper_A_En_c), .\control_reg[7] (control_reg_adj_1066[7]), 
            .n12211(n12211), .Stepper_A_Step_c(Stepper_A_Step_c), .limit_c_3(limit_c_3), 
            .n8654(n8653[7]), .n31410(n31410), .n8402(n8402), .n8368(n8368), 
            .n16843(n16843)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(625[25] 638[45])
    LUT4 Select_4229_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n31502), .C(read_value_adj_1107[28]), 
         .D(n33385), .Z(n8_adj_909)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4229_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    
endmodule
//
// Verilog Description of module ExpansionGPIO
//

module ExpansionGPIO (read_value, debug_c_c, n2870, n29221, n13948, 
            n31512, \databus[0] , \read_size[0] , n27680, prev_select, 
            \select[5] , expansion1_c_9, n31436, n56, expansion2_c_10, 
            expansion3_c_11, \databus[1] , \databus[2] , \databus[3] , 
            \register[0][4] , \databus[4] , \register[0][5] , \databus[5] , 
            \databus[6] , \databus[7] , n16013, \register[1][4] , \register[1][5] , 
            n12369, n31407, \register_addr[0] , n24146, n11008, n11007) /* synthesis syn_module_defined=1 */ ;
    output [7:0]read_value;
    input debug_c_c;
    input n2870;
    input n29221;
    input n13948;
    input n31512;
    input \databus[0] ;
    output \read_size[0] ;
    input n27680;
    output prev_select;
    input \select[5] ;
    output expansion1_c_9;
    input n31436;
    input n56;
    output expansion2_c_10;
    output expansion3_c_11;
    input \databus[1] ;
    input \databus[2] ;
    input \databus[3] ;
    output \register[0][4] ;
    input \databus[4] ;
    output \register[0][5] ;
    input \databus[5] ;
    input \databus[6] ;
    input \databus[7] ;
    input n16013;
    output \register[1][4] ;
    output \register[1][5] ;
    input n12369;
    input n31407;
    input \register_addr[0] ;
    input n24146;
    output n11008;
    output n11007;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [7:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(17[12:20])
    wire [7:0]n7637;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(17[12:20])
    wire [7:0]n7662;
    
    FD1P3AX read_value_i0_i4 (.D(n29221), .SP(n2870), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i4.GSR = "ENABLED";
    FD1P3IX register_0___i1 (.D(\databus[0] ), .SP(n13948), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i1.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n27680), .SP(n2870), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1S3AX prev_select_145 (.D(\select[5] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam prev_select_145.GSR = "ENABLED";
    LUT4 mux_2028_i2_4_lut (.A(expansion1_c_9), .B(\register[0] [1]), .C(n31436), 
         .D(n56), .Z(n7637[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2028_i2_4_lut.init = 16'ha0ac;
    LUT4 mux_2028_i3_4_lut (.A(expansion2_c_10), .B(\register[0] [2]), .C(n31436), 
         .D(n56), .Z(n7637[2])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2028_i3_4_lut.init = 16'ha0ac;
    LUT4 mux_2028_i4_4_lut (.A(expansion3_c_11), .B(\register[0] [3]), .C(n31436), 
         .D(n56), .Z(n7637[3])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2028_i4_4_lut.init = 16'ha0ac;
    FD1P3IX register_0___i2 (.D(\databus[1] ), .SP(n13948), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i2.GSR = "ENABLED";
    FD1P3IX register_0___i3 (.D(\databus[2] ), .SP(n13948), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i3.GSR = "ENABLED";
    FD1P3IX register_0___i4 (.D(\databus[3] ), .SP(n13948), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i4.GSR = "ENABLED";
    FD1P3IX register_0___i5 (.D(\databus[4] ), .SP(n13948), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[0][4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i5.GSR = "ENABLED";
    FD1P3IX register_0___i6 (.D(\databus[5] ), .SP(n13948), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[0][5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i6.GSR = "ENABLED";
    FD1P3IX register_0___i7 (.D(\databus[6] ), .SP(n13948), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i7.GSR = "ENABLED";
    FD1P3IX register_0___i8 (.D(\databus[7] ), .SP(n13948), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i8.GSR = "ENABLED";
    FD1P3IX register_0___i9 (.D(\databus[0] ), .SP(n16013), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i9.GSR = "ENABLED";
    FD1P3IX register_0___i10 (.D(\databus[1] ), .SP(n16013), .CD(n31512), 
            .CK(debug_c_c), .Q(expansion1_c_9)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i10.GSR = "ENABLED";
    FD1P3IX register_0___i11 (.D(\databus[2] ), .SP(n16013), .CD(n31512), 
            .CK(debug_c_c), .Q(expansion2_c_10)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i11.GSR = "ENABLED";
    FD1P3IX register_0___i12 (.D(\databus[3] ), .SP(n16013), .CD(n31512), 
            .CK(debug_c_c), .Q(expansion3_c_11)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i12.GSR = "ENABLED";
    FD1P3IX register_0___i13 (.D(\databus[4] ), .SP(n16013), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[1][4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i13.GSR = "ENABLED";
    FD1P3IX register_0___i14 (.D(\databus[5] ), .SP(n16013), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[1][5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i14.GSR = "ENABLED";
    FD1P3IX register_0___i15 (.D(\databus[6] ), .SP(n16013), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i15.GSR = "ENABLED";
    FD1P3IX register_0___i16 (.D(\databus[7] ), .SP(n12369), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i16.GSR = "ENABLED";
    FD1P3AX read_value_i0_i1 (.D(n7637[1]), .SP(n2870), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i1.GSR = "ENABLED";
    FD1P3AX read_value_i0_i2 (.D(n7637[2]), .SP(n2870), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i2.GSR = "ENABLED";
    FD1P3AX read_value_i0_i3 (.D(n7637[3]), .SP(n2870), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i3.GSR = "ENABLED";
    FD1P3AX read_value_i0_i5 (.D(n31407), .SP(n2870), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i5.GSR = "ENABLED";
    LUT4 mux_2029_Mux_7_i1_3_lut (.A(\register[0] [7]), .B(\register[1] [7]), 
         .C(\register_addr[0] ), .Z(n7662[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2029_Mux_7_i1_3_lut.init = 16'hcaca;
    LUT4 mux_2029_Mux_6_i1_3_lut (.A(\register[0] [6]), .B(\register[1] [6]), 
         .C(\register_addr[0] ), .Z(n7662[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2029_Mux_6_i1_3_lut.init = 16'hcaca;
    FD1P3IX read_value_i0_i7 (.D(n7662[7]), .SP(n2870), .CD(n24146), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i7.GSR = "ENABLED";
    FD1P3IX read_value_i0_i6 (.D(n7662[6]), .SP(n2870), .CD(n24146), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i6.GSR = "ENABLED";
    FD1P3IX read_value_i0_i0 (.D(n7662[0]), .SP(n2870), .CD(n24146), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i0.GSR = "ENABLED";
    LUT4 mux_2029_Mux_0_i1_3_lut (.A(\register[0] [0]), .B(\register[1] [0]), 
         .C(\register_addr[0] ), .Z(n7662[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2029_Mux_0_i1_3_lut.init = 16'hcaca;
    LUT4 Select_4215_i3_4_lut (.A(\register[1][4] ), .B(\register[0][5] ), 
         .C(\register[0][4] ), .D(\register[1][5] ), .Z(n11008)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam Select_4215_i3_4_lut.init = 16'heca0;
    LUT4 i22469_2_lut (.A(\register[0][5] ), .B(\register[0][4] ), .Z(n11007)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i22469_2_lut.init = 16'h1111;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0100000) 
//

module \ArmPeripheral(axis_haddr=8'b0100000)  (read_value, debug_c_c, n2847, 
            GND_net, VCC_net, Stepper_Z_nFault_c, n31512, \read_size[0] , 
            n27753, Stepper_Z_M0_c_0, n31420, databus, limit_latched, 
            prev_limit_latched, n9305, prev_select, n31483, \read_size[2] , 
            n29301, \register_addr[1] , \register_addr[5] , n31497, 
            rw, \select[4] , n52, \read_size[0]_adj_312 , n5, prev_select_adj_313, 
            n31422, \steps_reg[7] , n31601, n31556, n31591, n31596, 
            \register_addr[4] , n29271, n31464, Stepper_Z_M1_c_1, \register_addr[0] , 
            n29235, n31504, \read_size[2]_adj_314 , n9, Stepper_Z_M2_c_2, 
            n14523, n610, n608, Stepper_Z_Dir_c, Stepper_Z_En_c, n11209, 
            n14547, \register_addr[3] , \register_addr[2] , n31541, 
            n6, n4007, Stepper_Z_Step_c, limit_c_2, n11, n31411, 
            n16842, n8264, n8298) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    input n2847;
    input GND_net;
    input VCC_net;
    input Stepper_Z_nFault_c;
    input n31512;
    output \read_size[0] ;
    input n27753;
    output Stepper_Z_M0_c_0;
    input n31420;
    input [31:0]databus;
    output limit_latched;
    output prev_limit_latched;
    input n9305;
    output prev_select;
    input n31483;
    output \read_size[2] ;
    input n29301;
    input \register_addr[1] ;
    input \register_addr[5] ;
    input n31497;
    input rw;
    input \select[4] ;
    output n52;
    input \read_size[0]_adj_312 ;
    output n5;
    input prev_select_adj_313;
    output n31422;
    output \steps_reg[7] ;
    input n31601;
    input n31556;
    output n31591;
    input n31596;
    input \register_addr[4] ;
    output n29271;
    output n31464;
    output Stepper_Z_M1_c_1;
    input \register_addr[0] ;
    input n29235;
    input n31504;
    input \read_size[2]_adj_314 ;
    output n9;
    output Stepper_Z_M2_c_2;
    input n14523;
    input n610;
    input n608;
    output Stepper_Z_Dir_c;
    output Stepper_Z_En_c;
    input n11209;
    input n14547;
    input \register_addr[3] ;
    input \register_addr[2] ;
    output n31541;
    output n6;
    input n4007;
    output Stepper_Z_Step_c;
    input limit_c_2;
    input n11;
    input n31411;
    input n16842;
    output n8264;
    output n8298;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n31617, n26846;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n224;
    
    wire n26847, n26845, n26844, n26843, fault_latched;
    wire [31:0]n4008;
    
    wire prev_step_clk, step_clk, n182;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n31616, n31615, n26842, n26841, n26840, n26839, n26838, 
        n26837, n26836, n19911;
    wire [31:0]n100;
    
    wire n21, n17, n19, n19931, n29770, n29719, n27422;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n49, n62_adj_595, n58_adj_596, n50, n41, n60_adj_597, n54_adj_598, 
        n42_adj_599, n52_adj_600, n38_adj_601, n56_adj_602, n46_adj_603, 
        n29717, n29718, n27421, n29768, n29769, n19929;
    wire [7:0]n8644;
    
    wire int_step;
    wire [31:0]n7057;
    
    wire n10, n31418, n26851, n26850, n26849, n26848;
    
    FD1P3AX read_value__i0 (.D(n31617), .SP(n2847), .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26846), .COUT(n26847), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26845), .COUT(n26846), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26844), .COUT(n26845), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26843), .COUT(n26844), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    IFS1P3DX fault_latched_178 (.D(Stepper_Z_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n4008[0]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n27753), .SP(n2847), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3IX control_reg_i1 (.D(databus[0]), .SP(n31420), .CD(n31512), 
            .CK(debug_c_c), .Q(Stepper_Z_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i0 (.D(databus[0]), .SP(n9305), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n31483), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n29301), .SP(n2847), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n4008[31]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n4008[30]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n4008[29]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n4008[28]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n4008[27]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n4008[26]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n4008[25]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    LUT4 n30930_bdd_4_lut_then_3_lut (.A(steps_reg[0]), .B(limit_latched), 
         .C(\register_addr[1] ), .Z(n31616)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n30930_bdd_4_lut_then_3_lut.init = 16'hacac;
    LUT4 n30930_bdd_4_lut_else_3_lut (.A(Stepper_Z_M0_c_0), .B(div_factor_reg[0]), 
         .C(\register_addr[1] ), .Z(n31615)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30930_bdd_4_lut_else_3_lut.init = 16'hcaca;
    LUT4 i20_2_lut_3_lut_4_lut (.A(\register_addr[5] ), .B(n31497), .C(rw), 
         .D(\select[4] ), .Z(n52)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i20_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\register_addr[5] ), .B(n31497), .C(\read_size[0]_adj_312 ), 
         .D(\select[4] ), .Z(n5)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_rep_278_3_lut_4_lut (.A(\register_addr[5] ), .B(n31497), 
         .C(prev_select_adj_313), .D(\select[4] ), .Z(n31422)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_rep_278_3_lut_4_lut.init = 16'h0400;
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26842), .COUT(n26843), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26841), .COUT(n26842), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26840), .COUT(n26841), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(\steps_reg[7] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26839), .COUT(n26840), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26838), .COUT(n26839), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26837), .COUT(n26838), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26836), .COUT(n26837), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(step_clk), .C1(n19911), .D1(prev_step_clk), 
          .COUT(n26836), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n100[26]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n21), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n100[20]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n17), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n19), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n19931), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n29770), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n29719), .SP(n2847), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i2_3_lut (.A(n27422), .B(n31601), .C(control_reg[7]), .Z(n19911)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i2_3_lut.init = 16'h2020;
    LUT4 i31_4_lut (.A(n49), .B(n62_adj_595), .C(n58_adj_596), .D(n50), 
         .Z(n27422)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[15]), .B(steps_reg[23]), .C(steps_reg[21]), 
         .D(steps_reg[31]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60_adj_597), .C(n54_adj_598), .D(n42_adj_599), 
         .Z(n62_adj_595)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_504 (.A(n31556), .B(n31591), .C(n31596), 
         .D(\register_addr[4] ), .Z(n29271)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(83[9:13])
    defparam i1_2_lut_3_lut_4_lut_adj_504.init = 16'h0100;
    LUT4 i1_2_lut_rep_320_3_lut_4_lut (.A(n31556), .B(n31591), .C(n31596), 
         .D(\register_addr[4] ), .Z(n31464)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(83[9:13])
    defparam i1_2_lut_rep_320_3_lut_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[27]), .B(n52_adj_600), .C(n38_adj_601), 
         .D(steps_reg[20]), .Z(n58_adj_596)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[29]), .B(steps_reg[14]), .C(steps_reg[30]), 
         .D(steps_reg[19]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[16]), .B(steps_reg[24]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[8]), .B(n56_adj_602), .C(n46_adj_603), 
         .D(steps_reg[0]), .Z(n60_adj_597)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[9]), .B(steps_reg[17]), .C(steps_reg[12]), 
         .D(steps_reg[2]), .Z(n54_adj_598)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[25]), .B(steps_reg[26]), .Z(n42_adj_599)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[6]), .B(steps_reg[4]), .C(steps_reg[10]), 
         .D(steps_reg[3]), .Z(n56_adj_602)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[22]), .B(steps_reg[5]), .Z(n46_adj_603)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[13]), .B(steps_reg[18]), .C(steps_reg[28]), 
         .D(steps_reg[1]), .Z(n52_adj_600)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[11]), .B(\steps_reg[7] ), .Z(n38_adj_601)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i22157_3_lut (.A(Stepper_Z_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n29717)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22157_3_lut.init = 16'hcaca;
    LUT4 i22158_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n29718)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22158_3_lut.init = 16'hcaca;
    LUT4 i14897_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14897_4_lut.init = 16'hc088;
    LUT4 i14898_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14898_4_lut.init = 16'hc088;
    LUT4 i14899_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14899_4_lut.init = 16'hc088;
    LUT4 i1_4_lut (.A(\register_addr[1] ), .B(div_factor_reg[27]), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_4_lut.init = 16'ha088;
    LUT4 i14900_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n100[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14900_4_lut.init = 16'hc088;
    LUT4 i14901_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14901_4_lut.init = 16'hc088;
    LUT4 i14902_4_lut (.A(div_factor_reg[24]), .B(\register_addr[1] ), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14902_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_505 (.A(\register_addr[1] ), .B(div_factor_reg[23]), 
         .C(steps_reg[23]), .D(\register_addr[0] ), .Z(n21)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_4_lut_adj_505.init = 16'ha088;
    LUT4 i14903_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14903_4_lut.init = 16'hc088;
    LUT4 i14904_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14904_4_lut.init = 16'hc088;
    LUT4 i14905_4_lut (.A(div_factor_reg[20]), .B(\register_addr[1] ), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n100[20])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14905_4_lut.init = 16'hc088;
    LUT4 i14906_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14906_4_lut.init = 16'hc088;
    LUT4 i14907_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14907_4_lut.init = 16'hc088;
    LUT4 i14908_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14908_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_506 (.A(\register_addr[1] ), .B(div_factor_reg[16]), 
         .C(steps_reg[16]), .D(\register_addr[0] ), .Z(n17)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_4_lut_adj_506.init = 16'ha088;
    LUT4 i1_4_lut_adj_507 (.A(\register_addr[1] ), .B(div_factor_reg[15]), 
         .C(steps_reg[15]), .D(\register_addr[0] ), .Z(n19)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_4_lut_adj_507.init = 16'ha088;
    LUT4 i14909_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14909_4_lut.init = 16'hc088;
    LUT4 i14910_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14910_4_lut.init = 16'hc088;
    LUT4 i14911_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14911_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_508 (.A(\select[4] ), .B(n29235), .C(n31504), .D(\read_size[2]_adj_314 ), 
         .Z(n9)) /* synthesis lut_function=(A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut_adj_508.init = 16'h8a88;
    LUT4 i14912_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14912_4_lut.init = 16'hc088;
    LUT4 i14913_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14913_4_lut.init = 16'hc088;
    LUT4 i14914_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14914_4_lut.init = 16'hc088;
    LUT4 i14915_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14915_4_lut.init = 16'hc088;
    LUT4 i2_4_lut_4_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), 
         .C(steps_reg[31]), .D(div_factor_reg[31]), .Z(n27421)) /* synthesis lut_function=(A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i2_4_lut_4_lut.init = 16'ha280;
    FD1S3IX steps_reg__i24 (.D(n4008[24]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n4008[23]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n4008[22]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n4008[21]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n4008[20]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n4008[19]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n4008[18]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n4008[17]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n4008[16]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n4008[15]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n4008[14]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n4008[13]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n4008[12]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n4008[11]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n4008[10]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n4008[9]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n4008[8]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n4008[7]), .CK(debug_c_c), .CD(n31512), 
            .Q(\steps_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n4008[6]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n4008[5]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n4008[4]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n4008[3]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n4008[2]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n4008[1]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    PFUMX i22210 (.BLUT(n29768), .ALUT(n29769), .C0(\register_addr[0] ), 
          .Z(n29770));
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n31420), .PD(n31512), 
            .CK(debug_c_c), .Q(Stepper_Z_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n14523), .CK(debug_c_c), .Q(Stepper_Z_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n31420), .PD(n31512), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n14523), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n31420), .PD(n31512), 
            .CK(debug_c_c), .Q(Stepper_Z_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n31420), .PD(n31512), 
            .CK(debug_c_c), .Q(Stepper_Z_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n31420), .CD(n11209), 
            .CK(debug_c_c), .Q(control_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n14547), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n14547), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n9305), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n9305), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n9305), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n9305), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n9305), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n9305), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n9305), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n9305), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n9305), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n9305), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n9305), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n9305), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n9305), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n9305), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n9305), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n9305), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 i13172_3_lut (.A(control_reg[7]), .B(div_factor_reg[7]), .C(\register_addr[1] ), 
         .Z(n19929)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i13172_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_447 (.A(\register_addr[1] ), .B(\register_addr[0] ), 
         .Z(n31591)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(83[9:13])
    defparam i1_2_lut_rep_447.init = 16'heeee;
    LUT4 i2_2_lut_rep_397_3_lut_4_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), 
         .C(\register_addr[3] ), .D(\register_addr[2] ), .Z(n31541)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(83[9:13])
    defparam i2_2_lut_rep_397_3_lut_4_lut.init = 16'hfffe;
    LUT4 equal_67_i8_1_lut_2_lut_3_lut_4_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), 
         .C(\register_addr[3] ), .D(\register_addr[2] ), .Z(n6)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(83[9:13])
    defparam equal_67_i8_1_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    PFUMX i22159 (.BLUT(n29717), .ALUT(n29718), .C0(\register_addr[1] ), 
          .Z(n29719));
    LUT4 mux_1576_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n4007), 
         .Z(n4008[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n4007), 
         .Z(n4008[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n4007), 
         .Z(n4008[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n4007), 
         .Z(n4008[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n4007), 
         .Z(n4008[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n4007), 
         .Z(n4008[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n4007), 
         .Z(n4008[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n4007), 
         .Z(n4008[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n4007), 
         .Z(n4008[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n4007), 
         .Z(n4008[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n4007), 
         .Z(n4008[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n4007), 
         .Z(n4008[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n4007), 
         .Z(n4008[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n4007), 
         .Z(n4008[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n4007), 
         .Z(n4008[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n4007), .Z(n4008[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n4007), .Z(n4008[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n4007), .Z(n4008[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n4007), .Z(n4008[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n4007), .Z(n4008[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n4007), .Z(n4008[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n4007), .Z(n4008[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n4007), .Z(n4008[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n4007), .Z(n4008[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i2_3_lut.init = 16'hcaca;
    LUT4 i14927_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n8644[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14927_2_lut.init = 16'h2222;
    FD1P3AX read_value__i31 (.D(n27421), .SP(n2847), .CK(debug_c_c), .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_Z_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 mux_1976_i4_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), .C(\register_addr[0] ), 
         .Z(n7057[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1976_i4_3_lut.init = 16'hcaca;
    FD1P3AX int_step_182 (.D(n31418), .SP(n10), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 mux_1576_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n4007), .Z(n4008[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i1_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n14547), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n14547), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n14547), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n14547), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n14547), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n14547), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n14547), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n14547), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n14547), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n14547), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n14547), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n14547), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n14547), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    LUT4 i14926_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n8644[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14926_2_lut.init = 16'h2222;
    LUT4 i118_1_lut (.A(limit_c_2), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 mux_1976_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n7057[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1976_i5_3_lut.init = 16'hcaca;
    LUT4 i14925_2_lut (.A(Stepper_Z_Dir_c), .B(\register_addr[0] ), .Z(n8644[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14925_2_lut.init = 16'h2222;
    LUT4 i22208_3_lut (.A(Stepper_Z_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n29768)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22208_3_lut.init = 16'hcaca;
    LUT4 mux_1976_i6_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), .C(\register_addr[0] ), 
         .Z(n7057[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1976_i6_3_lut.init = 16'hcaca;
    LUT4 i22209_3_lut (.A(n19911), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n29769)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22209_3_lut.init = 16'hcaca;
    LUT4 i14924_2_lut (.A(Stepper_Z_En_c), .B(\register_addr[0] ), .Z(n8644[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14924_2_lut.init = 16'h2222;
    LUT4 mux_1976_i7_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n7057[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1976_i7_3_lut.init = 16'hcaca;
    PFUMX i13174 (.BLUT(n19929), .ALUT(n11), .C0(\register_addr[0] ), 
          .Z(n19931));
    LUT4 mux_1576_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n4007), 
         .Z(n4008[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n4007), 
         .Z(n4008[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n4007), 
         .Z(n4008[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n4007), 
         .Z(n4008[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n4007), 
         .Z(n4008[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n4007), 
         .Z(n4008[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1576_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n4007), 
         .Z(n4008[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1576_i26_3_lut.init = 16'hcaca;
    PFUMX mux_1980_i4 (.BLUT(n8644[3]), .ALUT(n7057[3]), .C0(\register_addr[1] ), 
          .Z(n100[3]));
    PFUMX mux_1980_i5 (.BLUT(n8644[4]), .ALUT(n7057[4]), .C0(\register_addr[1] ), 
          .Z(n100[4]));
    PFUMX mux_1980_i6 (.BLUT(n8644[5]), .ALUT(n7057[5]), .C0(\register_addr[1] ), 
          .Z(n100[5]));
    PFUMX mux_1980_i7 (.BLUT(n8644[6]), .ALUT(n7057[6]), .C0(\register_addr[1] ), 
          .Z(n100[6]));
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26851), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26850), .COUT(n26851), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26849), .COUT(n26850), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    PFUMX i22984 (.BLUT(n31615), .ALUT(n31616), .C0(\register_addr[0] ), 
          .Z(n31617));
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26848), .COUT(n26849), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26847), .COUT(n26848), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    ClockDivider step_clk_gen (.prev_step_clk(prev_step_clk), .n19911(n19911), 
            .step_clk(step_clk), .n31418(n31418), .n31512(n31512), .n10(n10), 
            .debug_c_c(debug_c_c), .n31411(n31411), .GND_net(GND_net), 
            .n16842(n16842), .div_factor_reg({div_factor_reg}), .n8264(n8264), 
            .n8298(n8298)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider
//

module ClockDivider (prev_step_clk, n19911, step_clk, n31418, n31512, 
            n10, debug_c_c, n31411, GND_net, n16842, div_factor_reg, 
            n8264, n8298) /* synthesis syn_module_defined=1 */ ;
    input prev_step_clk;
    input n19911;
    output step_clk;
    output n31418;
    input n31512;
    output n10;
    input debug_c_c;
    input n31411;
    input GND_net;
    input n16842;
    input [31:0]div_factor_reg;
    output n8264;
    output n8298;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n8229;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n26603, n26602;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n26601, n26600, n26599, n26598, n26597, n26596, n26595, 
        n26594, n26593, n26592, n26591, n26590, n26589, n26588, 
        n26787;
    wire [31:0]n40;
    
    wire n26786, n26587, n26586, n26585, n26584, n26923, n26922, 
        n26785, n26583, n26582, n26784, n26783, n26921, n26581, 
        n26920, n26919, n26918, n26782, n26917, n26916, n26915, 
        n26914, n26781, n26580, n26780, n26913, n26579, n26912, 
        n26578, n26911, n26577, n26779, n26778, n26910, n26777, 
        n26909, n26908, n26776, n26775, n26576, n26575, n26774, 
        n26574, n26773, n26573, n26572, n26772, n26571, n26570, 
        n26569, n26568, n26567, n26566, n26565, n26564, n26563, 
        n26562, n26561, n26560, n26559, n26558, n26557, n26556;
    
    LUT4 i2_3_lut_rep_274 (.A(prev_step_clk), .B(n19911), .C(step_clk), 
         .Z(n31418)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam i2_3_lut_rep_274.init = 16'h4040;
    LUT4 i1_4_lut_4_lut (.A(prev_step_clk), .B(n19911), .C(step_clk), 
         .D(n31512), .Z(n10)) /* synthesis lut_function=(!(A (C+(D))+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam i1_4_lut_4_lut.init = 16'h004a;
    FD1S3IX clk_o_22 (.D(n8229), .CK(debug_c_c), .CD(n31512), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    FD1S3IX count_2676__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i0.GSR = "ENABLED";
    CCU2D sub_2074_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26603), .S1(n8229));
    defparam sub_2074_add_2_33.INIT0 = 16'h5555;
    defparam sub_2074_add_2_33.INIT1 = 16'h0000;
    defparam sub_2074_add_2_33.INJECT1_0 = "NO";
    defparam sub_2074_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26602), .COUT(n26603));
    defparam sub_2074_add_2_31.INIT0 = 16'h5999;
    defparam sub_2074_add_2_31.INIT1 = 16'h5999;
    defparam sub_2074_add_2_31.INJECT1_0 = "NO";
    defparam sub_2074_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26601), .COUT(n26602));
    defparam sub_2074_add_2_29.INIT0 = 16'h5999;
    defparam sub_2074_add_2_29.INIT1 = 16'h5999;
    defparam sub_2074_add_2_29.INJECT1_0 = "NO";
    defparam sub_2074_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26600), .COUT(n26601));
    defparam sub_2074_add_2_27.INIT0 = 16'h5999;
    defparam sub_2074_add_2_27.INIT1 = 16'h5999;
    defparam sub_2074_add_2_27.INJECT1_0 = "NO";
    defparam sub_2074_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26599), .COUT(n26600));
    defparam sub_2074_add_2_25.INIT0 = 16'h5999;
    defparam sub_2074_add_2_25.INIT1 = 16'h5999;
    defparam sub_2074_add_2_25.INJECT1_0 = "NO";
    defparam sub_2074_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26598), .COUT(n26599));
    defparam sub_2074_add_2_23.INIT0 = 16'h5999;
    defparam sub_2074_add_2_23.INIT1 = 16'h5999;
    defparam sub_2074_add_2_23.INJECT1_0 = "NO";
    defparam sub_2074_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26597), .COUT(n26598));
    defparam sub_2074_add_2_21.INIT0 = 16'h5999;
    defparam sub_2074_add_2_21.INIT1 = 16'h5999;
    defparam sub_2074_add_2_21.INJECT1_0 = "NO";
    defparam sub_2074_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26596), .COUT(n26597));
    defparam sub_2074_add_2_19.INIT0 = 16'h5999;
    defparam sub_2074_add_2_19.INIT1 = 16'h5999;
    defparam sub_2074_add_2_19.INJECT1_0 = "NO";
    defparam sub_2074_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26595), .COUT(n26596));
    defparam sub_2074_add_2_17.INIT0 = 16'h5999;
    defparam sub_2074_add_2_17.INIT1 = 16'h5999;
    defparam sub_2074_add_2_17.INJECT1_0 = "NO";
    defparam sub_2074_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26594), .COUT(n26595));
    defparam sub_2074_add_2_15.INIT0 = 16'h5999;
    defparam sub_2074_add_2_15.INIT1 = 16'h5999;
    defparam sub_2074_add_2_15.INJECT1_0 = "NO";
    defparam sub_2074_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26593), .COUT(n26594));
    defparam sub_2074_add_2_13.INIT0 = 16'h5999;
    defparam sub_2074_add_2_13.INIT1 = 16'h5999;
    defparam sub_2074_add_2_13.INJECT1_0 = "NO";
    defparam sub_2074_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26592), .COUT(n26593));
    defparam sub_2074_add_2_11.INIT0 = 16'h5999;
    defparam sub_2074_add_2_11.INIT1 = 16'h5999;
    defparam sub_2074_add_2_11.INJECT1_0 = "NO";
    defparam sub_2074_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26591), .COUT(n26592));
    defparam sub_2074_add_2_9.INIT0 = 16'h5999;
    defparam sub_2074_add_2_9.INIT1 = 16'h5999;
    defparam sub_2074_add_2_9.INJECT1_0 = "NO";
    defparam sub_2074_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26590), .COUT(n26591));
    defparam sub_2074_add_2_7.INIT0 = 16'h5999;
    defparam sub_2074_add_2_7.INIT1 = 16'h5999;
    defparam sub_2074_add_2_7.INJECT1_0 = "NO";
    defparam sub_2074_add_2_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_2074_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26589), .COUT(n26590));
    defparam sub_2074_add_2_5.INIT0 = 16'h5999;
    defparam sub_2074_add_2_5.INIT1 = 16'h5999;
    defparam sub_2074_add_2_5.INJECT1_0 = "NO";
    defparam sub_2074_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26588), .COUT(n26589));
    defparam sub_2074_add_2_3.INIT0 = 16'h5999;
    defparam sub_2074_add_2_3.INIT1 = 16'h5999;
    defparam sub_2074_add_2_3.INJECT1_0 = "NO";
    defparam sub_2074_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26787), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26786), .COUT(n26787), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26588));
    defparam sub_2074_add_2_1.INIT0 = 16'h0000;
    defparam sub_2074_add_2_1.INIT1 = 16'h5999;
    defparam sub_2074_add_2_1.INJECT1_0 = "NO";
    defparam sub_2074_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26587), .S1(n8264));
    defparam sub_2076_add_2_33.INIT0 = 16'h5999;
    defparam sub_2076_add_2_33.INIT1 = 16'h0000;
    defparam sub_2076_add_2_33.INJECT1_0 = "NO";
    defparam sub_2076_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26586), .COUT(n26587));
    defparam sub_2076_add_2_31.INIT0 = 16'h5999;
    defparam sub_2076_add_2_31.INIT1 = 16'h5999;
    defparam sub_2076_add_2_31.INJECT1_0 = "NO";
    defparam sub_2076_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26585), .COUT(n26586));
    defparam sub_2076_add_2_29.INIT0 = 16'h5999;
    defparam sub_2076_add_2_29.INIT1 = 16'h5999;
    defparam sub_2076_add_2_29.INJECT1_0 = "NO";
    defparam sub_2076_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26584), .COUT(n26585));
    defparam sub_2076_add_2_27.INIT0 = 16'h5999;
    defparam sub_2076_add_2_27.INIT1 = 16'h5999;
    defparam sub_2076_add_2_27.INJECT1_0 = "NO";
    defparam sub_2076_add_2_27.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26923), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_33.INIT1 = 16'h0000;
    defparam count_2676_add_4_33.INJECT1_0 = "NO";
    defparam count_2676_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26922), .COUT(n26923), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_31.INJECT1_0 = "NO";
    defparam count_2676_add_4_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26785), .COUT(n26786), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26583), .COUT(n26584));
    defparam sub_2076_add_2_25.INIT0 = 16'h5999;
    defparam sub_2076_add_2_25.INIT1 = 16'h5999;
    defparam sub_2076_add_2_25.INJECT1_0 = "NO";
    defparam sub_2076_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26582), .COUT(n26583));
    defparam sub_2076_add_2_23.INIT0 = 16'h5999;
    defparam sub_2076_add_2_23.INIT1 = 16'h5999;
    defparam sub_2076_add_2_23.INJECT1_0 = "NO";
    defparam sub_2076_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26784), .COUT(n26785), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26783), .COUT(n26784), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26921), .COUT(n26922), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_29.INJECT1_0 = "NO";
    defparam count_2676_add_4_29.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26581), .COUT(n26582));
    defparam sub_2076_add_2_21.INIT0 = 16'h5999;
    defparam sub_2076_add_2_21.INIT1 = 16'h5999;
    defparam sub_2076_add_2_21.INJECT1_0 = "NO";
    defparam sub_2076_add_2_21.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26920), .COUT(n26921), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_27.INJECT1_0 = "NO";
    defparam count_2676_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26919), .COUT(n26920), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_25.INJECT1_0 = "NO";
    defparam count_2676_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26918), .COUT(n26919), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_23.INJECT1_0 = "NO";
    defparam count_2676_add_4_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26782), .COUT(n26783), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26917), .COUT(n26918), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_21.INJECT1_0 = "NO";
    defparam count_2676_add_4_21.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    CCU2D count_2676_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26916), .COUT(n26917), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_19.INJECT1_0 = "NO";
    defparam count_2676_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26915), .COUT(n26916), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_17.INJECT1_0 = "NO";
    defparam count_2676_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26914), .COUT(n26915), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_15.INJECT1_0 = "NO";
    defparam count_2676_add_4_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26781), .COUT(n26782), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    CCU2D sub_2076_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26580), .COUT(n26581));
    defparam sub_2076_add_2_19.INIT0 = 16'h5999;
    defparam sub_2076_add_2_19.INIT1 = 16'h5999;
    defparam sub_2076_add_2_19.INJECT1_0 = "NO";
    defparam sub_2076_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26780), .COUT(n26781), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26913), .COUT(n26914), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_13.INJECT1_0 = "NO";
    defparam count_2676_add_4_13.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26579), .COUT(n26580));
    defparam sub_2076_add_2_17.INIT0 = 16'h5999;
    defparam sub_2076_add_2_17.INIT1 = 16'h5999;
    defparam sub_2076_add_2_17.INJECT1_0 = "NO";
    defparam sub_2076_add_2_17.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    CCU2D count_2676_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26912), .COUT(n26913), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_11.INJECT1_0 = "NO";
    defparam count_2676_add_4_11.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26578), .COUT(n26579));
    defparam sub_2076_add_2_15.INIT0 = 16'h5999;
    defparam sub_2076_add_2_15.INIT1 = 16'h5999;
    defparam sub_2076_add_2_15.INJECT1_0 = "NO";
    defparam sub_2076_add_2_15.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26911), .COUT(n26912), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_9.INJECT1_0 = "NO";
    defparam count_2676_add_4_9.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26577), .COUT(n26578));
    defparam sub_2076_add_2_13.INIT0 = 16'h5999;
    defparam sub_2076_add_2_13.INIT1 = 16'h5999;
    defparam sub_2076_add_2_13.INJECT1_0 = "NO";
    defparam sub_2076_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26779), .COUT(n26780), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26778), .COUT(n26779), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26910), .COUT(n26911), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_7.INJECT1_0 = "NO";
    defparam count_2676_add_4_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26777), .COUT(n26778), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26909), .COUT(n26910), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_5.INJECT1_0 = "NO";
    defparam count_2676_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26908), .COUT(n26909), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2676_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2676_add_4_3.INJECT1_0 = "NO";
    defparam count_2676_add_4_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26776), .COUT(n26777), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D count_2676_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26908), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676_add_4_1.INIT0 = 16'hF000;
    defparam count_2676_add_4_1.INIT1 = 16'h0555;
    defparam count_2676_add_4_1.INJECT1_0 = "NO";
    defparam count_2676_add_4_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26775), .COUT(n26776), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26576), .COUT(n26577));
    defparam sub_2076_add_2_11.INIT0 = 16'h5999;
    defparam sub_2076_add_2_11.INIT1 = 16'h5999;
    defparam sub_2076_add_2_11.INJECT1_0 = "NO";
    defparam sub_2076_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26575), .COUT(n26576));
    defparam sub_2076_add_2_9.INIT0 = 16'h5999;
    defparam sub_2076_add_2_9.INIT1 = 16'h5999;
    defparam sub_2076_add_2_9.INJECT1_0 = "NO";
    defparam sub_2076_add_2_9.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26774), .COUT(n26775), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31411), .CD(n16842), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31411), .PD(n16842), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_2076_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26574), .COUT(n26575));
    defparam sub_2076_add_2_7.INIT0 = 16'h5999;
    defparam sub_2076_add_2_7.INIT1 = 16'h5999;
    defparam sub_2076_add_2_7.INJECT1_0 = "NO";
    defparam sub_2076_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26773), .COUT(n26774), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    FD1S3IX count_2676__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i1.GSR = "ENABLED";
    CCU2D sub_2076_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26573), .COUT(n26574));
    defparam sub_2076_add_2_5.INIT0 = 16'h5999;
    defparam sub_2076_add_2_5.INIT1 = 16'h5999;
    defparam sub_2076_add_2_5.INJECT1_0 = "NO";
    defparam sub_2076_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26572), .COUT(n26573));
    defparam sub_2076_add_2_3.INIT0 = 16'h5999;
    defparam sub_2076_add_2_3.INIT1 = 16'h5999;
    defparam sub_2076_add_2_3.INJECT1_0 = "NO";
    defparam sub_2076_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2076_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n26572));
    defparam sub_2076_add_2_1.INIT0 = 16'h0000;
    defparam sub_2076_add_2_1.INIT1 = 16'h5999;
    defparam sub_2076_add_2_1.INJECT1_0 = "NO";
    defparam sub_2076_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26772), .COUT(n26773), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26571), .S1(n8298));
    defparam sub_2077_add_2_33.INIT0 = 16'hf555;
    defparam sub_2077_add_2_33.INIT1 = 16'h0000;
    defparam sub_2077_add_2_33.INJECT1_0 = "NO";
    defparam sub_2077_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26772), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26570), .COUT(n26571));
    defparam sub_2077_add_2_31.INIT0 = 16'hf555;
    defparam sub_2077_add_2_31.INIT1 = 16'hf555;
    defparam sub_2077_add_2_31.INJECT1_0 = "NO";
    defparam sub_2077_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26569), .COUT(n26570));
    defparam sub_2077_add_2_29.INIT0 = 16'hf555;
    defparam sub_2077_add_2_29.INIT1 = 16'hf555;
    defparam sub_2077_add_2_29.INJECT1_0 = "NO";
    defparam sub_2077_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26568), .COUT(n26569));
    defparam sub_2077_add_2_27.INIT0 = 16'hf555;
    defparam sub_2077_add_2_27.INIT1 = 16'hf555;
    defparam sub_2077_add_2_27.INJECT1_0 = "NO";
    defparam sub_2077_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26567), .COUT(n26568));
    defparam sub_2077_add_2_25.INIT0 = 16'hf555;
    defparam sub_2077_add_2_25.INIT1 = 16'hf555;
    defparam sub_2077_add_2_25.INJECT1_0 = "NO";
    defparam sub_2077_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26566), .COUT(n26567));
    defparam sub_2077_add_2_23.INIT0 = 16'hf555;
    defparam sub_2077_add_2_23.INIT1 = 16'hf555;
    defparam sub_2077_add_2_23.INJECT1_0 = "NO";
    defparam sub_2077_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26565), .COUT(n26566));
    defparam sub_2077_add_2_21.INIT0 = 16'hf555;
    defparam sub_2077_add_2_21.INIT1 = 16'hf555;
    defparam sub_2077_add_2_21.INJECT1_0 = "NO";
    defparam sub_2077_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26564), .COUT(n26565));
    defparam sub_2077_add_2_19.INIT0 = 16'hf555;
    defparam sub_2077_add_2_19.INIT1 = 16'hf555;
    defparam sub_2077_add_2_19.INJECT1_0 = "NO";
    defparam sub_2077_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26563), .COUT(n26564));
    defparam sub_2077_add_2_17.INIT0 = 16'hf555;
    defparam sub_2077_add_2_17.INIT1 = 16'hf555;
    defparam sub_2077_add_2_17.INJECT1_0 = "NO";
    defparam sub_2077_add_2_17.INJECT1_1 = "NO";
    FD1S3IX count_2676__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i2.GSR = "ENABLED";
    FD1S3IX count_2676__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i3.GSR = "ENABLED";
    FD1S3IX count_2676__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i4.GSR = "ENABLED";
    FD1S3IX count_2676__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i5.GSR = "ENABLED";
    FD1S3IX count_2676__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i6.GSR = "ENABLED";
    FD1S3IX count_2676__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i7.GSR = "ENABLED";
    FD1S3IX count_2676__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i8.GSR = "ENABLED";
    FD1S3IX count_2676__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i9.GSR = "ENABLED";
    FD1S3IX count_2676__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i10.GSR = "ENABLED";
    FD1S3IX count_2676__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i11.GSR = "ENABLED";
    FD1S3IX count_2676__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i12.GSR = "ENABLED";
    FD1S3IX count_2676__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i13.GSR = "ENABLED";
    FD1S3IX count_2676__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i14.GSR = "ENABLED";
    FD1S3IX count_2676__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i15.GSR = "ENABLED";
    FD1S3IX count_2676__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i16.GSR = "ENABLED";
    FD1S3IX count_2676__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i17.GSR = "ENABLED";
    FD1S3IX count_2676__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i18.GSR = "ENABLED";
    FD1S3IX count_2676__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i19.GSR = "ENABLED";
    FD1S3IX count_2676__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i20.GSR = "ENABLED";
    FD1S3IX count_2676__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i21.GSR = "ENABLED";
    FD1S3IX count_2676__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i22.GSR = "ENABLED";
    FD1S3IX count_2676__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i23.GSR = "ENABLED";
    FD1S3IX count_2676__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i24.GSR = "ENABLED";
    FD1S3IX count_2676__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i25.GSR = "ENABLED";
    FD1S3IX count_2676__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i26.GSR = "ENABLED";
    FD1S3IX count_2676__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i27.GSR = "ENABLED";
    FD1S3IX count_2676__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i28.GSR = "ENABLED";
    FD1S3IX count_2676__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i29.GSR = "ENABLED";
    FD1S3IX count_2676__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i30.GSR = "ENABLED";
    FD1S3IX count_2676__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31411), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2676__i31.GSR = "ENABLED";
    CCU2D sub_2077_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26562), .COUT(n26563));
    defparam sub_2077_add_2_15.INIT0 = 16'hf555;
    defparam sub_2077_add_2_15.INIT1 = 16'hf555;
    defparam sub_2077_add_2_15.INJECT1_0 = "NO";
    defparam sub_2077_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26561), .COUT(n26562));
    defparam sub_2077_add_2_13.INIT0 = 16'hf555;
    defparam sub_2077_add_2_13.INIT1 = 16'hf555;
    defparam sub_2077_add_2_13.INJECT1_0 = "NO";
    defparam sub_2077_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26560), .COUT(n26561));
    defparam sub_2077_add_2_11.INIT0 = 16'hf555;
    defparam sub_2077_add_2_11.INIT1 = 16'hf555;
    defparam sub_2077_add_2_11.INJECT1_0 = "NO";
    defparam sub_2077_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26559), .COUT(n26560));
    defparam sub_2077_add_2_9.INIT0 = 16'hf555;
    defparam sub_2077_add_2_9.INIT1 = 16'hf555;
    defparam sub_2077_add_2_9.INJECT1_0 = "NO";
    defparam sub_2077_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26558), .COUT(n26559));
    defparam sub_2077_add_2_7.INIT0 = 16'hf555;
    defparam sub_2077_add_2_7.INIT1 = 16'hf555;
    defparam sub_2077_add_2_7.INJECT1_0 = "NO";
    defparam sub_2077_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26557), .COUT(n26558));
    defparam sub_2077_add_2_5.INIT0 = 16'hf555;
    defparam sub_2077_add_2_5.INIT1 = 16'hf555;
    defparam sub_2077_add_2_5.INJECT1_0 = "NO";
    defparam sub_2077_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26556), .COUT(n26557));
    defparam sub_2077_add_2_3.INIT0 = 16'hf555;
    defparam sub_2077_add_2_3.INIT1 = 16'hf555;
    defparam sub_2077_add_2_3.INJECT1_0 = "NO";
    defparam sub_2077_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2077_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n26556));
    defparam sub_2077_add_2_1.INIT0 = 16'h0000;
    defparam sub_2077_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2077_add_2_1.INJECT1_0 = "NO";
    defparam sub_2077_add_2_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b010000) 
//

module \ArmPeripheral(axis_haddr=8'b010000)  (debug_c_c, VCC_net, GND_net, 
            Stepper_Y_nFault_c, n31512, n4095, \read_size[0] , n14651, 
            n27752, Stepper_Y_M0_c_0, databus, prev_step_clk, step_clk, 
            limit_latched, prev_limit_latched, n9301, prev_select, n31446, 
            n29271, n29492, Stepper_Y_M1_c_1, \register_addr[0] , \div_factor_reg[9] , 
            \div_factor_reg[6] , \div_factor_reg[5] , \div_factor_reg[4] , 
            \div_factor_reg[3] , \control_reg[7] , n12149, Stepper_Y_En_c, 
            Stepper_Y_Dir_c, \control_reg[4] , \control_reg[3] , Stepper_Y_M2_c_2, 
            \read_size[2] , n29200, \steps_reg[9] , \steps_reg[6] , 
            \steps_reg[5] , \steps_reg[4] , \steps_reg[3] , read_value, 
            n9548, \register_addr[1] , n29113, limit_c_1, int_step, 
            n22, n31419, n29114, n21214, n21222, n28827, n6808, 
            n32, n27484, n224, n8636, n8194, n31408, n16841, n8160) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input VCC_net;
    input GND_net;
    input Stepper_Y_nFault_c;
    input n31512;
    input [31:0]n4095;
    output \read_size[0] ;
    input n14651;
    input n27752;
    output Stepper_Y_M0_c_0;
    input [31:0]databus;
    output prev_step_clk;
    output step_clk;
    output limit_latched;
    output prev_limit_latched;
    input n9301;
    output prev_select;
    input n31446;
    input n29271;
    input n29492;
    output Stepper_Y_M1_c_1;
    input \register_addr[0] ;
    output \div_factor_reg[9] ;
    output \div_factor_reg[6] ;
    output \div_factor_reg[5] ;
    output \div_factor_reg[4] ;
    output \div_factor_reg[3] ;
    output \control_reg[7] ;
    input n12149;
    output Stepper_Y_En_c;
    output Stepper_Y_Dir_c;
    output \control_reg[4] ;
    output \control_reg[3] ;
    output Stepper_Y_M2_c_2;
    output \read_size[2] ;
    input n29200;
    output \steps_reg[9] ;
    output \steps_reg[6] ;
    output \steps_reg[5] ;
    output \steps_reg[4] ;
    output \steps_reg[3] ;
    output [31:0]read_value;
    input n9548;
    input \register_addr[1] ;
    input n29113;
    input limit_c_1;
    output int_step;
    input n22;
    input n31419;
    input n29114;
    input n21214;
    input n21222;
    input n28827;
    input n6808;
    input n32;
    output n27484;
    output [31:0]n224;
    input n8636;
    output n8194;
    input n31408;
    input n16841;
    output n8160;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire fault_latched;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire n13924, n182;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n29714, n29715, n29741, n29742, n29743;
    wire [31:0]n100;
    
    wire n29687, n29688, n29689, n29716;
    wire [31:0]n6743;
    
    wire n29133, n29121, n29134, n29135, n29136, n29132, n29131, 
        n29130, n29129, n29126, n29128, n29127, n29125, n29124, 
        n29123, n29122, n29115, n29119, n29117, n29120, n29118, 
        n29116;
    wire [31:0]n6779;
    
    wire n49, n62, n58, n50, n41, n60, n54, n42, n52, n38, 
        n56, n46, n26867, n26866, n26865, n26864, n26863, n26862, 
        n26861, n26860, n26859, n26858, n26857, n26856, n26855, 
        n26854, n26853, n26852;
    
    IFS1P3DX fault_latched_178 (.D(Stepper_Y_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n4095[0]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n27752), .SP(n14651), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3IX control_reg_i1 (.D(databus[0]), .SP(n13924), .CD(n31512), 
            .CK(debug_c_c), .Q(Stepper_Y_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i0 (.D(databus[0]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n31446), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(n31446), .B(prev_select), .C(n29271), 
         .D(n29492), .Z(n13924)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i22154_3_lut (.A(Stepper_Y_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n29714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22154_3_lut.init = 16'hcaca;
    LUT4 i22155_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n29715)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22155_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n9301), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n9301), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n9301), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n9301), .PD(n31512), 
            .CK(debug_c_c), .Q(\div_factor_reg[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n9301), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n9301), .PD(n31512), 
            .CK(debug_c_c), .Q(\div_factor_reg[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n9301), .PD(n31512), 
            .CK(debug_c_c), .Q(\div_factor_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(\div_factor_reg[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(\div_factor_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n9301), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n13924), .CD(n12149), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n13924), .PD(n31512), 
            .CK(debug_c_c), .Q(Stepper_Y_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n13924), .PD(n31512), 
            .CK(debug_c_c), .Q(Stepper_Y_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n13924), .CD(n31512), 
            .CK(debug_c_c), .Q(\control_reg[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n13924), .PD(n31512), 
            .CK(debug_c_c), .Q(\control_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n13924), .CD(n31512), 
            .CK(debug_c_c), .Q(Stepper_Y_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n13924), .PD(n31512), 
            .CK(debug_c_c), .Q(Stepper_Y_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    PFUMX i22183 (.BLUT(n29741), .ALUT(n29742), .C0(\register_addr[0] ), 
          .Z(n29743));
    FD1P3AX read_size__i2 (.D(n29200), .SP(n14651), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n4095[31]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n4095[30]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n4095[29]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n4095[28]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n4095[27]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n4095[26]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n4095[25]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n4095[24]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n4095[23]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n4095[22]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n4095[21]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n4095[20]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n4095[19]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n4095[18]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n4095[17]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n4095[16]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n4095[15]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n4095[14]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n4095[13]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n4095[12]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n4095[11]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n4095[10]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n4095[9]), .CK(debug_c_c), .CD(n31512), 
            .Q(\steps_reg[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n4095[8]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n4095[7]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n4095[6]), .CK(debug_c_c), .CD(n31512), 
            .Q(\steps_reg[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n4095[5]), .CK(debug_c_c), .CD(n31512), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n4095[4]), .CK(debug_c_c), .CD(n31512), 
            .Q(\steps_reg[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n4095[3]), .CK(debug_c_c), .CD(n31512), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n4095[2]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n4095[1]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n14651), .CD(n9548), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    PFUMX i22129 (.BLUT(n29687), .ALUT(n29688), .C0(\register_addr[1] ), 
          .Z(n29689));
    PFUMX i22156 (.BLUT(n29714), .ALUT(n29715), .C0(\register_addr[1] ), 
          .Z(n29716));
    LUT4 i22127_3_lut (.A(Stepper_Y_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n29687)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22127_3_lut.init = 16'hcaca;
    LUT4 i22128_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n29688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22128_3_lut.init = 16'hcaca;
    LUT4 mux_1950_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n6743[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1950_i8_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i30 (.D(n29133), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n29121), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n29134), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n29135), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n29136), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n29132), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29131), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29130), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29129), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29126), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29128), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n29127), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29125), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29124), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29123), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29122), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(div_factor_reg[30]), .B(n29113), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n29133)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i118_1_lut (.A(limit_c_1), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_483 (.A(div_factor_reg[29]), .B(n29113), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n29121)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_483.init = 16'hc088;
    FD1P3AX int_step_182 (.D(n31419), .SP(n22), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29115), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29119), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29117), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29120), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29118), .SP(n14651), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29114), .SP(n14651), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29116), .SP(n14651), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6779[7]), .SP(n14651), .CD(n9548), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n21214), .SP(n14651), .CD(n9548), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n21222), .SP(n14651), .CD(n9548), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n28827), .SP(n14651), .CD(n9548), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6808), .SP(n14651), .CD(n9548), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n29743), .SP(n14651), .CD(n9548), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n29716), .SP(n14651), .CD(n9548), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_484 (.A(div_factor_reg[28]), .B(n29113), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n29134)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_484.init = 16'hc088;
    LUT4 i1_4_lut_adj_485 (.A(div_factor_reg[27]), .B(n29113), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n29135)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_485.init = 16'hc088;
    LUT4 i1_4_lut_adj_486 (.A(div_factor_reg[26]), .B(n29113), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n29136)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_486.init = 16'hc088;
    LUT4 i1_4_lut_adj_487 (.A(div_factor_reg[25]), .B(n29113), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n29132)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_487.init = 16'hc088;
    LUT4 i1_4_lut_adj_488 (.A(div_factor_reg[24]), .B(n29113), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n29131)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_488.init = 16'hc088;
    LUT4 i1_4_lut_adj_489 (.A(div_factor_reg[23]), .B(n29113), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n29130)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_489.init = 16'hc088;
    LUT4 i1_4_lut_adj_490 (.A(div_factor_reg[22]), .B(n29113), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n29129)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_490.init = 16'hc088;
    LUT4 i22181_3_lut (.A(Stepper_Y_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n29741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22181_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i0 (.D(n29689), .SP(n14651), .CD(n9548), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i22182_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n29742)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22182_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_491 (.A(div_factor_reg[21]), .B(n29113), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n29126)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_491.init = 16'hc088;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n27484)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[0]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_492 (.A(div_factor_reg[20]), .B(n29113), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n29128)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_492.init = 16'hc088;
    LUT4 i1_4_lut_adj_493 (.A(div_factor_reg[19]), .B(n29113), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n29127)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_493.init = 16'hc088;
    LUT4 i1_4_lut_adj_494 (.A(div_factor_reg[18]), .B(n29113), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n29125)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_494.init = 16'hc088;
    LUT4 i1_4_lut_adj_495 (.A(div_factor_reg[17]), .B(n29113), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n29124)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_495.init = 16'hc088;
    LUT4 i1_4_lut_adj_496 (.A(div_factor_reg[16]), .B(n29113), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n29123)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_496.init = 16'hc088;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_497 (.A(div_factor_reg[15]), .B(n29113), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n29122)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_497.init = 16'hc088;
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52), .C(n38), .D(steps_reg[18]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[7]), .B(\steps_reg[5] ), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[26]), .B(n56), .C(n46), .D(steps_reg[29]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[24]), .B(\steps_reg[4] ), .C(steps_reg[1]), 
         .D(steps_reg[25]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[10]), .B(steps_reg[22]), .C(steps_reg[20]), 
         .D(\steps_reg[6] ), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(\steps_reg[9] ), .B(\steps_reg[3] ), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[28]), .C(steps_reg[13]), 
         .D(steps_reg[30]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[2]), .B(steps_reg[8]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_498 (.A(div_factor_reg[14]), .B(n29113), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n29115)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_498.init = 16'hc088;
    LUT4 i1_4_lut_adj_499 (.A(div_factor_reg[13]), .B(n29113), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n29119)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_499.init = 16'hc088;
    LUT4 i1_4_lut_adj_500 (.A(div_factor_reg[12]), .B(n29113), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n29117)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_500.init = 16'hc088;
    LUT4 i1_4_lut_adj_501 (.A(div_factor_reg[11]), .B(n29113), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n29120)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_501.init = 16'hc088;
    LUT4 i1_4_lut_adj_502 (.A(div_factor_reg[10]), .B(n29113), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n29118)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_502.init = 16'hc088;
    LUT4 i1_4_lut_adj_503 (.A(div_factor_reg[8]), .B(n29113), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n29116)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_503.init = 16'hc088;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26867), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26866), .COUT(n26867), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26865), .COUT(n26866), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26864), .COUT(n26865), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26863), .COUT(n26864), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26862), .COUT(n26863), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26861), .COUT(n26862), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26860), .COUT(n26861), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26859), .COUT(n26860), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26858), .COUT(n26859), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26857), .COUT(n26858), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(\steps_reg[9] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26856), .COUT(n26857), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    PFUMX mux_1954_i8 (.BLUT(n8636), .ALUT(n6743[7]), .C0(\register_addr[1] ), 
          .Z(n6779[7]));
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26855), .COUT(n26856), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    LUT4 i14928_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14928_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26854), .COUT(n26855), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[4] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26853), .COUT(n26854), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26852), .COUT(n26853), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n26852), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    ClockDivider_U7 step_clk_gen (.GND_net(GND_net), .step_clk(step_clk), 
            .debug_c_c(debug_c_c), .n31512(n31512), .div_factor_reg({div_factor_reg[31:10], 
            \div_factor_reg[9] , div_factor_reg[8:7], \div_factor_reg[6] , 
            \div_factor_reg[5] , \div_factor_reg[4] , \div_factor_reg[3] , 
            div_factor_reg[2:0]}), .n8194(n8194), .n31408(n31408), .n16841(n16841), 
            .n8160(n8160)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U7
//

module ClockDivider_U7 (GND_net, step_clk, debug_c_c, n31512, div_factor_reg, 
            n8194, n31408, n16841, n8160) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output step_clk;
    input debug_c_c;
    input n31512;
    input [31:0]div_factor_reg;
    output n8194;
    input n31408;
    input n16841;
    output n8160;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26629;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n40;
    
    wire n26630, n26628, n26627, n26626, n26625, n26624, n26623, 
        n26622, n8125, n26621, n26620, n26619, n26618, n26617, 
        n26616, n26615, n26614, n26613, n26612, n26611, n26610, 
        n26803;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n26609, n26802;
    wire [31:0]n134;
    
    wire n26801, n26800, n26799, n26798, n26797, n26608, n26796, 
        n26795, n26607, n26606, n26794, n26605, n26604, n26793, 
        n26792, n26791, n26790, n26789, n26788, n26651, n26650, 
        n26649, n26648, n26647, n26646, n26645, n26644, n27035, 
        n26643, n27034, n27033, n27032, n27031, n27030, n27029, 
        n27028, n27027, n26642, n26641, n27026, n27025, n27024, 
        n26640, n27023, n26639, n27022, n27021, n27020, n26638, 
        n26637, n26636, n26635, n26634, n26633, n26632, n26631;
    
    CCU2D sub_2071_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26629), .COUT(n26630));
    defparam sub_2071_add_2_21.INIT0 = 16'h5999;
    defparam sub_2071_add_2_21.INIT1 = 16'h5999;
    defparam sub_2071_add_2_21.INJECT1_0 = "NO";
    defparam sub_2071_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26628), .COUT(n26629));
    defparam sub_2071_add_2_19.INIT0 = 16'h5999;
    defparam sub_2071_add_2_19.INIT1 = 16'h5999;
    defparam sub_2071_add_2_19.INJECT1_0 = "NO";
    defparam sub_2071_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26627), .COUT(n26628));
    defparam sub_2071_add_2_17.INIT0 = 16'h5999;
    defparam sub_2071_add_2_17.INIT1 = 16'h5999;
    defparam sub_2071_add_2_17.INJECT1_0 = "NO";
    defparam sub_2071_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26626), .COUT(n26627));
    defparam sub_2071_add_2_15.INIT0 = 16'h5999;
    defparam sub_2071_add_2_15.INIT1 = 16'h5999;
    defparam sub_2071_add_2_15.INJECT1_0 = "NO";
    defparam sub_2071_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26625), .COUT(n26626));
    defparam sub_2071_add_2_13.INIT0 = 16'h5999;
    defparam sub_2071_add_2_13.INIT1 = 16'h5999;
    defparam sub_2071_add_2_13.INJECT1_0 = "NO";
    defparam sub_2071_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26624), .COUT(n26625));
    defparam sub_2071_add_2_11.INIT0 = 16'h5999;
    defparam sub_2071_add_2_11.INIT1 = 16'h5999;
    defparam sub_2071_add_2_11.INJECT1_0 = "NO";
    defparam sub_2071_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26623), .COUT(n26624));
    defparam sub_2071_add_2_9.INIT0 = 16'h5999;
    defparam sub_2071_add_2_9.INIT1 = 16'h5999;
    defparam sub_2071_add_2_9.INJECT1_0 = "NO";
    defparam sub_2071_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26622), .COUT(n26623));
    defparam sub_2071_add_2_7.INIT0 = 16'h5999;
    defparam sub_2071_add_2_7.INIT1 = 16'h5999;
    defparam sub_2071_add_2_7.INJECT1_0 = "NO";
    defparam sub_2071_add_2_7.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n8125), .CK(debug_c_c), .CD(n31512), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2071_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26621), .COUT(n26622));
    defparam sub_2071_add_2_5.INIT0 = 16'h5999;
    defparam sub_2071_add_2_5.INIT1 = 16'h5999;
    defparam sub_2071_add_2_5.INJECT1_0 = "NO";
    defparam sub_2071_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26620), .COUT(n26621));
    defparam sub_2071_add_2_3.INIT0 = 16'h5999;
    defparam sub_2071_add_2_3.INIT1 = 16'h5999;
    defparam sub_2071_add_2_3.INJECT1_0 = "NO";
    defparam sub_2071_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n26620));
    defparam sub_2071_add_2_1.INIT0 = 16'h0000;
    defparam sub_2071_add_2_1.INIT1 = 16'h5999;
    defparam sub_2071_add_2_1.INJECT1_0 = "NO";
    defparam sub_2071_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26619), .S1(n8194));
    defparam sub_2072_add_2_33.INIT0 = 16'hf555;
    defparam sub_2072_add_2_33.INIT1 = 16'h0000;
    defparam sub_2072_add_2_33.INJECT1_0 = "NO";
    defparam sub_2072_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26618), .COUT(n26619));
    defparam sub_2072_add_2_31.INIT0 = 16'hf555;
    defparam sub_2072_add_2_31.INIT1 = 16'hf555;
    defparam sub_2072_add_2_31.INJECT1_0 = "NO";
    defparam sub_2072_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26617), .COUT(n26618));
    defparam sub_2072_add_2_29.INIT0 = 16'hf555;
    defparam sub_2072_add_2_29.INIT1 = 16'hf555;
    defparam sub_2072_add_2_29.INJECT1_0 = "NO";
    defparam sub_2072_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26616), .COUT(n26617));
    defparam sub_2072_add_2_27.INIT0 = 16'hf555;
    defparam sub_2072_add_2_27.INIT1 = 16'hf555;
    defparam sub_2072_add_2_27.INJECT1_0 = "NO";
    defparam sub_2072_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26615), .COUT(n26616));
    defparam sub_2072_add_2_25.INIT0 = 16'hf555;
    defparam sub_2072_add_2_25.INIT1 = 16'hf555;
    defparam sub_2072_add_2_25.INJECT1_0 = "NO";
    defparam sub_2072_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26614), .COUT(n26615));
    defparam sub_2072_add_2_23.INIT0 = 16'hf555;
    defparam sub_2072_add_2_23.INIT1 = 16'hf555;
    defparam sub_2072_add_2_23.INJECT1_0 = "NO";
    defparam sub_2072_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26613), .COUT(n26614));
    defparam sub_2072_add_2_21.INIT0 = 16'hf555;
    defparam sub_2072_add_2_21.INIT1 = 16'hf555;
    defparam sub_2072_add_2_21.INJECT1_0 = "NO";
    defparam sub_2072_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26612), .COUT(n26613));
    defparam sub_2072_add_2_19.INIT0 = 16'hf555;
    defparam sub_2072_add_2_19.INIT1 = 16'hf555;
    defparam sub_2072_add_2_19.INJECT1_0 = "NO";
    defparam sub_2072_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26611), .COUT(n26612));
    defparam sub_2072_add_2_17.INIT0 = 16'hf555;
    defparam sub_2072_add_2_17.INIT1 = 16'hf555;
    defparam sub_2072_add_2_17.INJECT1_0 = "NO";
    defparam sub_2072_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26610), .COUT(n26611));
    defparam sub_2072_add_2_15.INIT0 = 16'hf555;
    defparam sub_2072_add_2_15.INIT1 = 16'hf555;
    defparam sub_2072_add_2_15.INJECT1_0 = "NO";
    defparam sub_2072_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26803), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26609), .COUT(n26610));
    defparam sub_2072_add_2_13.INIT0 = 16'hf555;
    defparam sub_2072_add_2_13.INIT1 = 16'hf555;
    defparam sub_2072_add_2_13.INJECT1_0 = "NO";
    defparam sub_2072_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26802), .COUT(n26803), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    FD1S3IX count_2675__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i0.GSR = "ENABLED";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26801), .COUT(n26802), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26800), .COUT(n26801), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26799), .COUT(n26800), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26798), .COUT(n26799), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26797), .COUT(n26798), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26608), .COUT(n26609));
    defparam sub_2072_add_2_11.INIT0 = 16'hf555;
    defparam sub_2072_add_2_11.INIT1 = 16'hf555;
    defparam sub_2072_add_2_11.INJECT1_0 = "NO";
    defparam sub_2072_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26796), .COUT(n26797), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26795), .COUT(n26796), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26607), .COUT(n26608));
    defparam sub_2072_add_2_9.INIT0 = 16'hf555;
    defparam sub_2072_add_2_9.INIT1 = 16'hf555;
    defparam sub_2072_add_2_9.INJECT1_0 = "NO";
    defparam sub_2072_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26606), .COUT(n26607));
    defparam sub_2072_add_2_7.INIT0 = 16'hf555;
    defparam sub_2072_add_2_7.INIT1 = 16'hf555;
    defparam sub_2072_add_2_7.INJECT1_0 = "NO";
    defparam sub_2072_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26794), .COUT(n26795), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26605), .COUT(n26606));
    defparam sub_2072_add_2_5.INIT0 = 16'hf555;
    defparam sub_2072_add_2_5.INIT1 = 16'hf555;
    defparam sub_2072_add_2_5.INJECT1_0 = "NO";
    defparam sub_2072_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26604), .COUT(n26605));
    defparam sub_2072_add_2_3.INIT0 = 16'hf555;
    defparam sub_2072_add_2_3.INIT1 = 16'hf555;
    defparam sub_2072_add_2_3.INJECT1_0 = "NO";
    defparam sub_2072_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26793), .COUT(n26794), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n26604));
    defparam sub_2072_add_2_1.INIT0 = 16'h0000;
    defparam sub_2072_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2072_add_2_1.INJECT1_0 = "NO";
    defparam sub_2072_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26792), .COUT(n26793), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26791), .COUT(n26792), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26790), .COUT(n26791), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26789), .COUT(n26790), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26788), .COUT(n26789), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26788), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31408), .CD(n16841), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31408), .PD(n16841), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_2069_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26651), .S1(n8125));
    defparam sub_2069_add_2_33.INIT0 = 16'h5555;
    defparam sub_2069_add_2_33.INIT1 = 16'h0000;
    defparam sub_2069_add_2_33.INJECT1_0 = "NO";
    defparam sub_2069_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26650), .COUT(n26651));
    defparam sub_2069_add_2_31.INIT0 = 16'h5999;
    defparam sub_2069_add_2_31.INIT1 = 16'h5999;
    defparam sub_2069_add_2_31.INJECT1_0 = "NO";
    defparam sub_2069_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26649), .COUT(n26650));
    defparam sub_2069_add_2_29.INIT0 = 16'h5999;
    defparam sub_2069_add_2_29.INIT1 = 16'h5999;
    defparam sub_2069_add_2_29.INJECT1_0 = "NO";
    defparam sub_2069_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26648), .COUT(n26649));
    defparam sub_2069_add_2_27.INIT0 = 16'h5999;
    defparam sub_2069_add_2_27.INIT1 = 16'h5999;
    defparam sub_2069_add_2_27.INJECT1_0 = "NO";
    defparam sub_2069_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26647), .COUT(n26648));
    defparam sub_2069_add_2_25.INIT0 = 16'h5999;
    defparam sub_2069_add_2_25.INIT1 = 16'h5999;
    defparam sub_2069_add_2_25.INJECT1_0 = "NO";
    defparam sub_2069_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26646), .COUT(n26647));
    defparam sub_2069_add_2_23.INIT0 = 16'h5999;
    defparam sub_2069_add_2_23.INIT1 = 16'h5999;
    defparam sub_2069_add_2_23.INJECT1_0 = "NO";
    defparam sub_2069_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26645), .COUT(n26646));
    defparam sub_2069_add_2_21.INIT0 = 16'h5999;
    defparam sub_2069_add_2_21.INIT1 = 16'h5999;
    defparam sub_2069_add_2_21.INJECT1_0 = "NO";
    defparam sub_2069_add_2_21.INJECT1_1 = "NO";
    FD1S3IX count_2675__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i1.GSR = "ENABLED";
    FD1S3IX count_2675__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i2.GSR = "ENABLED";
    FD1S3IX count_2675__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i3.GSR = "ENABLED";
    FD1S3IX count_2675__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i4.GSR = "ENABLED";
    FD1S3IX count_2675__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i5.GSR = "ENABLED";
    FD1S3IX count_2675__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i6.GSR = "ENABLED";
    FD1S3IX count_2675__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i7.GSR = "ENABLED";
    FD1S3IX count_2675__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i8.GSR = "ENABLED";
    FD1S3IX count_2675__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i9.GSR = "ENABLED";
    FD1S3IX count_2675__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i10.GSR = "ENABLED";
    FD1S3IX count_2675__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i11.GSR = "ENABLED";
    FD1S3IX count_2675__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i12.GSR = "ENABLED";
    FD1S3IX count_2675__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i13.GSR = "ENABLED";
    FD1S3IX count_2675__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i14.GSR = "ENABLED";
    FD1S3IX count_2675__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i15.GSR = "ENABLED";
    FD1S3IX count_2675__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i16.GSR = "ENABLED";
    FD1S3IX count_2675__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i17.GSR = "ENABLED";
    FD1S3IX count_2675__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i18.GSR = "ENABLED";
    FD1S3IX count_2675__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i19.GSR = "ENABLED";
    FD1S3IX count_2675__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i20.GSR = "ENABLED";
    FD1S3IX count_2675__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i21.GSR = "ENABLED";
    FD1S3IX count_2675__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i22.GSR = "ENABLED";
    FD1S3IX count_2675__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i23.GSR = "ENABLED";
    FD1S3IX count_2675__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i24.GSR = "ENABLED";
    FD1S3IX count_2675__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i25.GSR = "ENABLED";
    FD1S3IX count_2675__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i26.GSR = "ENABLED";
    FD1S3IX count_2675__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i27.GSR = "ENABLED";
    FD1S3IX count_2675__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i28.GSR = "ENABLED";
    FD1S3IX count_2675__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i29.GSR = "ENABLED";
    FD1S3IX count_2675__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i30.GSR = "ENABLED";
    FD1S3IX count_2675__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31408), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675__i31.GSR = "ENABLED";
    CCU2D sub_2069_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26644), .COUT(n26645));
    defparam sub_2069_add_2_19.INIT0 = 16'h5999;
    defparam sub_2069_add_2_19.INIT1 = 16'h5999;
    defparam sub_2069_add_2_19.INJECT1_0 = "NO";
    defparam sub_2069_add_2_19.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27035), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_33.INIT1 = 16'h0000;
    defparam count_2675_add_4_33.INJECT1_0 = "NO";
    defparam count_2675_add_4_33.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26643), .COUT(n26644));
    defparam sub_2069_add_2_17.INIT0 = 16'h5999;
    defparam sub_2069_add_2_17.INIT1 = 16'h5999;
    defparam sub_2069_add_2_17.INJECT1_0 = "NO";
    defparam sub_2069_add_2_17.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27034), .COUT(n27035), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_31.INJECT1_0 = "NO";
    defparam count_2675_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27033), .COUT(n27034), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_29.INJECT1_0 = "NO";
    defparam count_2675_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27032), .COUT(n27033), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_27.INJECT1_0 = "NO";
    defparam count_2675_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27031), .COUT(n27032), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_25.INJECT1_0 = "NO";
    defparam count_2675_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27030), .COUT(n27031), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_23.INJECT1_0 = "NO";
    defparam count_2675_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27029), .COUT(n27030), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_21.INJECT1_0 = "NO";
    defparam count_2675_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27028), .COUT(n27029), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_19.INJECT1_0 = "NO";
    defparam count_2675_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27027), .COUT(n27028), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_17.INJECT1_0 = "NO";
    defparam count_2675_add_4_17.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26642), .COUT(n26643));
    defparam sub_2069_add_2_15.INIT0 = 16'h5999;
    defparam sub_2069_add_2_15.INIT1 = 16'h5999;
    defparam sub_2069_add_2_15.INJECT1_0 = "NO";
    defparam sub_2069_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26641), .COUT(n26642));
    defparam sub_2069_add_2_13.INIT0 = 16'h5999;
    defparam sub_2069_add_2_13.INIT1 = 16'h5999;
    defparam sub_2069_add_2_13.INJECT1_0 = "NO";
    defparam sub_2069_add_2_13.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27026), .COUT(n27027), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_15.INJECT1_0 = "NO";
    defparam count_2675_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27025), .COUT(n27026), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_13.INJECT1_0 = "NO";
    defparam count_2675_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27024), .COUT(n27025), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_11.INJECT1_0 = "NO";
    defparam count_2675_add_4_11.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26640), .COUT(n26641));
    defparam sub_2069_add_2_11.INIT0 = 16'h5999;
    defparam sub_2069_add_2_11.INIT1 = 16'h5999;
    defparam sub_2069_add_2_11.INJECT1_0 = "NO";
    defparam sub_2069_add_2_11.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27023), .COUT(n27024), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_9.INJECT1_0 = "NO";
    defparam count_2675_add_4_9.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26639), .COUT(n26640));
    defparam sub_2069_add_2_9.INIT0 = 16'h5999;
    defparam sub_2069_add_2_9.INIT1 = 16'h5999;
    defparam sub_2069_add_2_9.INJECT1_0 = "NO";
    defparam sub_2069_add_2_9.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27022), .COUT(n27023), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_7.INJECT1_0 = "NO";
    defparam count_2675_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27021), .COUT(n27022), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_5.INJECT1_0 = "NO";
    defparam count_2675_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27020), .COUT(n27021), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2675_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2675_add_4_3.INJECT1_0 = "NO";
    defparam count_2675_add_4_3.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26638), .COUT(n26639));
    defparam sub_2069_add_2_7.INIT0 = 16'h5999;
    defparam sub_2069_add_2_7.INIT1 = 16'h5999;
    defparam sub_2069_add_2_7.INJECT1_0 = "NO";
    defparam sub_2069_add_2_7.INJECT1_1 = "NO";
    CCU2D count_2675_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27020), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2675_add_4_1.INIT0 = 16'hF000;
    defparam count_2675_add_4_1.INIT1 = 16'h0555;
    defparam count_2675_add_4_1.INJECT1_0 = "NO";
    defparam count_2675_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26637), .COUT(n26638));
    defparam sub_2069_add_2_5.INIT0 = 16'h5999;
    defparam sub_2069_add_2_5.INIT1 = 16'h5999;
    defparam sub_2069_add_2_5.INJECT1_0 = "NO";
    defparam sub_2069_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26636), .COUT(n26637));
    defparam sub_2069_add_2_3.INIT0 = 16'h5999;
    defparam sub_2069_add_2_3.INIT1 = 16'h5999;
    defparam sub_2069_add_2_3.INJECT1_0 = "NO";
    defparam sub_2069_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26636));
    defparam sub_2069_add_2_1.INIT0 = 16'h0000;
    defparam sub_2069_add_2_1.INIT1 = 16'h5999;
    defparam sub_2069_add_2_1.INJECT1_0 = "NO";
    defparam sub_2069_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26635), .S1(n8160));
    defparam sub_2071_add_2_33.INIT0 = 16'h5999;
    defparam sub_2071_add_2_33.INIT1 = 16'h0000;
    defparam sub_2071_add_2_33.INJECT1_0 = "NO";
    defparam sub_2071_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26634), .COUT(n26635));
    defparam sub_2071_add_2_31.INIT0 = 16'h5999;
    defparam sub_2071_add_2_31.INIT1 = 16'h5999;
    defparam sub_2071_add_2_31.INJECT1_0 = "NO";
    defparam sub_2071_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26633), .COUT(n26634));
    defparam sub_2071_add_2_29.INIT0 = 16'h5999;
    defparam sub_2071_add_2_29.INIT1 = 16'h5999;
    defparam sub_2071_add_2_29.INJECT1_0 = "NO";
    defparam sub_2071_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26632), .COUT(n26633));
    defparam sub_2071_add_2_27.INIT0 = 16'h5999;
    defparam sub_2071_add_2_27.INIT1 = 16'h5999;
    defparam sub_2071_add_2_27.INJECT1_0 = "NO";
    defparam sub_2071_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26631), .COUT(n26632));
    defparam sub_2071_add_2_25.INIT0 = 16'h5999;
    defparam sub_2071_add_2_25.INIT1 = 16'h5999;
    defparam sub_2071_add_2_25.INJECT1_0 = "NO";
    defparam sub_2071_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2071_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26630), .COUT(n26631));
    defparam sub_2071_add_2_23.INIT0 = 16'h5999;
    defparam sub_2071_add_2_23.INIT1 = 16'h5999;
    defparam sub_2071_add_2_23.INJECT1_0 = "NO";
    defparam sub_2071_add_2_23.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module RCPeripheral
//

module RCPeripheral (n2, databus, \read_value[10] , n8, n31426, \register_addr[0] , 
            read_value, read_value_adj_308, n46, n52, databus_out, 
            rw, read_value_adj_309, \read_value[10]_adj_157 , n52_adj_158, 
            n31447, n2_adj_159, \read_value[9]_adj_160 , n8_adj_161, 
            \read_value[9]_adj_162 , n2_adj_163, \select[7] , n176, 
            \read_value[8]_adj_164 , n8_adj_165, \register_addr[1] , n2_adj_166, 
            \read_value[24]_adj_167 , n8_adj_168, \read_value[24]_adj_169 , 
            \read_value[8]_adj_170 , n2_adj_171, \read_value[7]_adj_172 , 
            \read_value[7]_adj_173 , n31444, n3, read_value_adj_310, 
            n64, n66, read_value_adj_311, \read_value[14]_adj_190 , 
            n2_adj_191, \read_value[6]_adj_192 , \read_value[6]_adj_193 , 
            n3_adj_194, n2_adj_195, \read_value[5]_adj_196 , \read_value[5]_adj_197 , 
            n33385, n3_adj_198, n2_adj_199, \read_value[4]_adj_200 , 
            \read_value[4]_adj_201 , n3_adj_202, n2_adj_203, \read_value[3]_adj_204 , 
            \read_value[3]_adj_205 , n2_adj_206, \read_value[22]_adj_207 , 
            n8_adj_208, n3_adj_209, n2_adj_210, \read_value[2]_adj_211 , 
            \read_value[2]_adj_212 , \read_value[22]_adj_213 , n3_adj_214, 
            n10, \read_value[1]_adj_215 , n3_adj_216, \read_value[1]_adj_217 , 
            n2_adj_218, \read_value[13]_adj_219 , n8_adj_220, n2_adj_221, 
            \read_value[13]_adj_222 , \read_value[23]_adj_223 , n8_adj_224, 
            n2_adj_225, n2_adj_226, \read_value[12]_adj_227 , n8_adj_228, 
            \read_value[23]_adj_229 , \read_value[12]_adj_230 , \read_value[21]_adj_231 , 
            n8_adj_232, read_size, \select[1] , n13, n31483, n9, 
            \read_size[0]_adj_233 , n18, \read_size[0]_adj_234 , \read_size[0]_adj_235 , 
            n31465, \select[2] , n14, n31474, n5, \read_size[0]_adj_236 , 
            \read_size[0]_adj_237 , n31445, \select[5] , \read_size[0]_adj_238 , 
            n2_adj_239, \read_value[11]_adj_240 , n8_adj_241, n6, \read_size[2]_adj_242 , 
            \reg_size[2] , \read_size[2]_adj_243 , n9_adj_244, \read_size[2]_adj_245 , 
            n31471, \read_value[11]_adj_246 , \read_value[21]_adj_247 , 
            n2_adj_248, \read_value[25]_adj_249 , n8_adj_250, \read_value[25]_adj_251 , 
            \register_addr[2] , n2_adj_252, n2_adj_253, \read_value[20]_adj_254 , 
            n8_adj_255, \read_value[16]_adj_256 , n8_adj_257, n31588, 
            \sendcount[1] , n13156, n31457, \read_value[20]_adj_258 , 
            n2_adj_259, n2_adj_260, \read_value[0]_adj_261 , \read_value[0]_adj_262 , 
            n3_adj_263, n2_adj_264, \read_value[26]_adj_265 , n8_adj_266, 
            \read_value[26]_adj_267 , \read_value[16]_adj_268 , n2_adj_269, 
            \read_value[19]_adj_270 , n8_adj_271, n29237, n2_adj_272, 
            \read_value[19]_adj_273 , n2_adj_274, \read_value[18]_adj_275 , 
            n8_adj_276, n2_adj_277, \read_value[31]_adj_278 , n8_adj_279, 
            \read_value[14]_adj_280 , n8_adj_281, \read_value[31]_adj_282 , 
            n2_adj_283, \read_value[30]_adj_284 , n8_adj_285, \read_value[18]_adj_286 , 
            \read_value[30]_adj_287 , n2_adj_288, \read_value[17]_adj_289 , 
            \read_value[29]_adj_290 , n8_adj_291, \read_value[29]_adj_292 , 
            n2_adj_293, n2_adj_294, \read_value[15]_adj_295 , n8_adj_296, 
            \read_value[28]_adj_297 , n8_adj_298, \read_value[17]_adj_299 , 
            n8_adj_300, \read_value[28]_adj_301 , n2_adj_302, \read_value[27]_adj_303 , 
            n8_adj_304, \read_value[15]_adj_305 , \read_value[27]_adj_306 , 
            GND_net, debug_c_c, n33387, rc_ch8_c, n29818, n33386, 
            n13957, n27564, n29784, rc_ch7_c, n33388, n27543, n29827, 
            rc_ch4_c, n27550, n29838, rc_ch3_c, n14500, n27541, 
            n29840, n29530, n29944, n14_adj_307, n29832, rc_ch2_c, 
            n31412, n14513, n29847, n27536, n31512, n14514, rc_ch1_c, 
            n29830, n27547, n29811) /* synthesis syn_module_defined=1 */ ;
    input n2;
    output [31:0]databus;
    input \read_value[10] ;
    input n8;
    input n31426;
    input \register_addr[0] ;
    input [31:0]read_value;
    input [31:0]read_value_adj_308;
    input n46;
    input n52;
    input [31:0]databus_out;
    input rw;
    input [31:0]read_value_adj_309;
    input \read_value[10]_adj_157 ;
    input n52_adj_158;
    input n31447;
    input n2_adj_159;
    input \read_value[9]_adj_160 ;
    input n8_adj_161;
    input \read_value[9]_adj_162 ;
    input n2_adj_163;
    input \select[7] ;
    input n176;
    input \read_value[8]_adj_164 ;
    input n8_adj_165;
    input \register_addr[1] ;
    input n2_adj_166;
    input \read_value[24]_adj_167 ;
    input n8_adj_168;
    input \read_value[24]_adj_169 ;
    input \read_value[8]_adj_170 ;
    input n2_adj_171;
    input \read_value[7]_adj_172 ;
    input \read_value[7]_adj_173 ;
    input n31444;
    input n3;
    input [7:0]read_value_adj_310;
    input n64;
    input n66;
    input [7:0]read_value_adj_311;
    input \read_value[14]_adj_190 ;
    input n2_adj_191;
    input \read_value[6]_adj_192 ;
    input \read_value[6]_adj_193 ;
    input n3_adj_194;
    input n2_adj_195;
    input \read_value[5]_adj_196 ;
    input \read_value[5]_adj_197 ;
    input n33385;
    input n3_adj_198;
    input n2_adj_199;
    input \read_value[4]_adj_200 ;
    input \read_value[4]_adj_201 ;
    input n3_adj_202;
    input n2_adj_203;
    input \read_value[3]_adj_204 ;
    input \read_value[3]_adj_205 ;
    input n2_adj_206;
    input \read_value[22]_adj_207 ;
    input n8_adj_208;
    input n3_adj_209;
    input n2_adj_210;
    input \read_value[2]_adj_211 ;
    input \read_value[2]_adj_212 ;
    input \read_value[22]_adj_213 ;
    input n3_adj_214;
    input n10;
    input \read_value[1]_adj_215 ;
    input n3_adj_216;
    input \read_value[1]_adj_217 ;
    input n2_adj_218;
    input \read_value[13]_adj_219 ;
    input n8_adj_220;
    input n2_adj_221;
    input \read_value[13]_adj_222 ;
    input \read_value[23]_adj_223 ;
    input n8_adj_224;
    input n2_adj_225;
    input n2_adj_226;
    input \read_value[12]_adj_227 ;
    input n8_adj_228;
    input \read_value[23]_adj_229 ;
    input \read_value[12]_adj_230 ;
    input \read_value[21]_adj_231 ;
    input n8_adj_232;
    input [2:0]read_size;
    input \select[1] ;
    output n13;
    input n31483;
    input n9;
    input \read_size[0]_adj_233 ;
    output n18;
    input \read_size[0]_adj_234 ;
    input \read_size[0]_adj_235 ;
    input n31465;
    input \select[2] ;
    output n14;
    input n31474;
    input n5;
    input \read_size[0]_adj_236 ;
    input \read_size[0]_adj_237 ;
    input n31445;
    input \select[5] ;
    input \read_size[0]_adj_238 ;
    input n2_adj_239;
    input \read_value[11]_adj_240 ;
    input n8_adj_241;
    input n6;
    input \read_size[2]_adj_242 ;
    output \reg_size[2] ;
    input \read_size[2]_adj_243 ;
    input n9_adj_244;
    input \read_size[2]_adj_245 ;
    input n31471;
    input \read_value[11]_adj_246 ;
    input \read_value[21]_adj_247 ;
    input n2_adj_248;
    input \read_value[25]_adj_249 ;
    input n8_adj_250;
    input \read_value[25]_adj_251 ;
    input \register_addr[2] ;
    input n2_adj_252;
    input n2_adj_253;
    input \read_value[20]_adj_254 ;
    input n8_adj_255;
    input \read_value[16]_adj_256 ;
    input n8_adj_257;
    output n31588;
    input \sendcount[1] ;
    output n13156;
    input n31457;
    input \read_value[20]_adj_258 ;
    input n2_adj_259;
    input n2_adj_260;
    input \read_value[0]_adj_261 ;
    input \read_value[0]_adj_262 ;
    input n3_adj_263;
    input n2_adj_264;
    input \read_value[26]_adj_265 ;
    input n8_adj_266;
    input \read_value[26]_adj_267 ;
    input \read_value[16]_adj_268 ;
    input n2_adj_269;
    input \read_value[19]_adj_270 ;
    input n8_adj_271;
    output n29237;
    input n2_adj_272;
    input \read_value[19]_adj_273 ;
    input n2_adj_274;
    input \read_value[18]_adj_275 ;
    input n8_adj_276;
    input n2_adj_277;
    input \read_value[31]_adj_278 ;
    input n8_adj_279;
    input \read_value[14]_adj_280 ;
    input n8_adj_281;
    input \read_value[31]_adj_282 ;
    input n2_adj_283;
    input \read_value[30]_adj_284 ;
    input n8_adj_285;
    input \read_value[18]_adj_286 ;
    input \read_value[30]_adj_287 ;
    input n2_adj_288;
    input \read_value[17]_adj_289 ;
    input \read_value[29]_adj_290 ;
    input n8_adj_291;
    input \read_value[29]_adj_292 ;
    input n2_adj_293;
    input n2_adj_294;
    input \read_value[15]_adj_295 ;
    input n8_adj_296;
    input \read_value[28]_adj_297 ;
    input n8_adj_298;
    input \read_value[17]_adj_299 ;
    input n8_adj_300;
    input \read_value[28]_adj_301 ;
    input n2_adj_302;
    input \read_value[27]_adj_303 ;
    input n8_adj_304;
    input \read_value[15]_adj_305 ;
    input \read_value[27]_adj_306 ;
    input GND_net;
    input debug_c_c;
    input n33387;
    input rc_ch8_c;
    output n29818;
    input n33386;
    input n13957;
    input n27564;
    output n29784;
    input rc_ch7_c;
    input n33388;
    input n27543;
    output n29827;
    input rc_ch4_c;
    input n27550;
    output n29838;
    input rc_ch3_c;
    input n14500;
    input n27541;
    output n29840;
    output n29530;
    output n29944;
    input n14_adj_307;
    output n29832;
    input rc_ch2_c;
    input n31412;
    input n14513;
    output n29847;
    input n27536;
    input n31512;
    input n14514;
    input rc_ch1_c;
    output n29830;
    input n27547;
    output n29811;
    
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(455[15:21])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n13_c, n11, n5_c, n10_c;
    wire [7:0]\register[6] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n30333, n13_adj_224, n11_adj_225, n5_adj_227, n10_adj_228, 
        n13_adj_234, n11_adj_235, n5_adj_237;
    wire [2:0]read_size_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(211[12:21])
    
    wire n10_adj_238, n30778, n30777, n30779;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n30337, n13_adj_240, n11_adj_241, n5_adj_243, n10_adj_244;
    wire [7:0]\register[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n30780, n1210, n30781, n15, n20, n7;
    wire [7:0]read_value_adj_588;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(210[12:22])
    
    wire n18_c, n12, n46_adj_257, n14_c, n5_adj_263, n10_adj_265, 
        n30816, n15_adj_266, n20_adj_267, n7_adj_269, n30817, n18_adj_272, 
        n12_adj_273, n14_adj_275, n30819, n15_adj_281, n20_adj_282, 
        n7_adj_284, n18_adj_287, n12_adj_288, n14_adj_290, n1225, 
        n30820, n15_adj_296, n20_adj_297, n7_adj_299, n18_adj_302, 
        n12_adj_303, n31157, n31155, n1240, n31158, n31154, n14_adj_305, 
        n15_adj_311, n20_adj_312, n7_adj_314, n18_adj_317, n12_adj_318, 
        n13_adj_319, n11_adj_320, n5_adj_322, n10_adj_323, n14_adj_328, 
        n30838, n30839, n15_adj_334, n20_adj_335, n7_adj_337, n30841, 
        n18_adj_340, n12_adj_341, n14_adj_345, n1195, n30842, n19, 
        n8_adj_351, n18_adj_352, n12_adj_353, n16, n14_adj_356, n13_adj_364, 
        n11_adj_365, n5_adj_367, n10_adj_368, n13_adj_370, n11_adj_371, 
        n5_adj_373, n10_adj_378, n30334, n13_adj_382, n11_adj_383, 
        n5_adj_385, n13_adj_386, n11_adj_387, n5_adj_389, n10_adj_390, 
        n10_adj_398, n16_adj_402, n12_adj_408, n13_adj_415, n11_adj_416, 
        n5_adj_418, n10_adj_419, n10_adj_423, n8_adj_425, n30888, 
        n30885, n30886, n1180, n30889, n31305, n31304, n31307, 
        n31308, n13_adj_433, n11_adj_434, n5_adj_436, n31317, n10_adj_437, 
        n31316, n31321, n31318, n31322, n31319, n31320, n1165, 
        n13_adj_443, n11_adj_444, n5_adj_446, n13_adj_447, n11_adj_448, 
        n5_adj_450, n10_adj_451, n10_adj_453, n31309, n31306, n31310, 
        n30891, n30844, n30783, n30339, n30822, n31160, n13_adj_461, 
        n11_adj_462, n15_adj_464, n20_adj_465, n7_adj_467, n18_adj_470, 
        n12_adj_471, n14_adj_473, n13_adj_475, n11_adj_476, n5_adj_478, 
        n10_adj_481, n30338, n30335, n31159, n31156, n13_adj_491, 
        n11_adj_492, n5_adj_494, n10_adj_495, n30336, n13_adj_499, 
        n11_adj_500, n5_adj_502, n30890, n30887, n13_adj_505, n11_adj_506, 
        n5_adj_508, n10_adj_509, n13_adj_513, n11_adj_514, n5_adj_516, 
        n10_adj_517, n5_adj_521, n13_adj_526, n11_adj_527, n5_adj_529, 
        n10_adj_530, n30843, n30840, n13_adj_538, n11_adj_539, n5_adj_541, 
        n10_adj_543, n10_adj_544, n13_adj_550, n11_adj_551, n5_adj_553, 
        n13_adj_556, n11_adj_557, n10_adj_559, n30821, n30818, n10_adj_563, 
        n13_adj_571, n11_adj_572, n5_adj_574, n10_adj_575, n30782;
    
    LUT4 i7_4_lut (.A(n13_c), .B(n11), .C(n2), .D(n5_c), .Z(databus[10])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i5_4_lut (.A(\read_value[10] ), .B(n10_c), .C(n8), .D(n31426), 
         .Z(n13_c)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_22611 (.A(\register[6] [5]), .B(\register_addr[0] ), 
         .Z(n30333)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22611.init = 16'h2222;
    LUT4 i3_4_lut (.A(read_value[10]), .B(read_value_adj_308[10]), .C(n46), 
         .D(n52), .Z(n11)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut.init = 16'heca0;
    LUT4 Select_4283_i5_2_lut (.A(databus_out[10]), .B(rw), .Z(n5_c)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4283_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut (.A(read_value_adj_309[10]), .B(\read_value[10]_adj_157 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut.init = 16'heca0;
    LUT4 i7_4_lut_adj_341 (.A(n13_adj_224), .B(n11_adj_225), .C(n2_adj_159), 
         .D(n5_adj_227), .Z(databus[9])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_341.init = 16'hfffe;
    LUT4 i5_4_lut_adj_342 (.A(\read_value[9]_adj_160 ), .B(n10_adj_228), 
         .C(n8_adj_161), .D(n31426), .Z(n13_adj_224)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_342.init = 16'hfefc;
    LUT4 i3_4_lut_adj_343 (.A(read_value[9]), .B(read_value_adj_308[9]), 
         .C(n46), .D(n52), .Z(n11_adj_225)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_343.init = 16'heca0;
    LUT4 Select_4286_i5_2_lut (.A(databus_out[9]), .B(rw), .Z(n5_adj_227)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4286_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_344 (.A(read_value_adj_309[9]), .B(\read_value[9]_adj_162 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_228)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_344.init = 16'heca0;
    LUT4 i7_4_lut_adj_345 (.A(n13_adj_234), .B(n11_adj_235), .C(n2_adj_163), 
         .D(n5_adj_237), .Z(databus[8])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_345.init = 16'hfffe;
    FD1S3AX read_size_i1 (.D(n176), .CK(\select[7] ), .Q(read_size_c[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_size_i1.GSR = "ENABLED";
    LUT4 i5_4_lut_adj_346 (.A(\read_value[8]_adj_164 ), .B(n10_adj_238), 
         .C(n8_adj_165), .D(n31426), .Z(n13_adj_234)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_346.init = 16'hfefc;
    PFUMX i22678 (.BLUT(n30778), .ALUT(n30777), .C0(\register_addr[1] ), 
          .Z(n30779));
    LUT4 \register_1[[5__bdd_2_lut_22782  (.A(\register[1] [5]), .B(\register_addr[0] ), 
         .Z(n30337)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[5__bdd_2_lut_22782 .init = 16'h8888;
    LUT4 i7_4_lut_adj_347 (.A(n13_adj_240), .B(n11_adj_241), .C(n2_adj_166), 
         .D(n5_adj_243), .Z(databus[24])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_347.init = 16'hfffe;
    LUT4 i5_4_lut_adj_348 (.A(\read_value[24]_adj_167 ), .B(n10_adj_244), 
         .C(n8_adj_168), .D(n31426), .Z(n13_adj_240)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_348.init = 16'hfefc;
    LUT4 register_addr_1__bdd_3_lut_22696 (.A(\register_addr[0] ), .B(\register[4] [3]), 
         .C(\register[5] [3]), .Z(n30778)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22696.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_22695 (.A(\register[6] [3]), .B(\register_addr[0] ), 
         .Z(n30777)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22695.init = 16'h2222;
    LUT4 i3_4_lut_adj_349 (.A(read_value[24]), .B(read_value_adj_308[24]), 
         .C(n46), .D(n52), .Z(n11_adj_241)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_349.init = 16'heca0;
    LUT4 n1210_bdd_3_lut_22680 (.A(\register[2] [3]), .B(\register[3] [3]), 
         .C(\register_addr[0] ), .Z(n30780)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1210_bdd_3_lut_22680.init = 16'hcaca;
    LUT4 Select_4241_i5_2_lut (.A(databus_out[24]), .B(rw), .Z(n5_adj_243)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4241_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_350 (.A(read_value_adj_309[24]), .B(\read_value[24]_adj_169 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_244)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_350.init = 16'heca0;
    LUT4 n1210_bdd_3_lut_22975 (.A(n1210), .B(\register_addr[0] ), .C(\register[1] [3]), 
         .Z(n30781)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1210_bdd_3_lut_22975.init = 16'he2e2;
    LUT4 i3_4_lut_adj_351 (.A(read_value[8]), .B(read_value_adj_308[8]), 
         .C(n46), .D(n52), .Z(n11_adj_235)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_351.init = 16'heca0;
    LUT4 Select_4289_i5_2_lut (.A(databus_out[8]), .B(rw), .Z(n5_adj_237)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4289_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_352 (.A(read_value_adj_309[8]), .B(\read_value[8]_adj_170 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_238)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_352.init = 16'heca0;
    LUT4 i10_4_lut (.A(n15), .B(n20), .C(n2_adj_171), .D(n7), .Z(databus[7])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i4_4_lut (.A(\read_value[7]_adj_172 ), .B(\read_value[7]_adj_173 ), 
         .C(n31447), .D(n31444), .Z(n15)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut.init = 16'heca0;
    LUT4 i9_4_lut (.A(read_value_adj_588[7]), .B(n18_c), .C(n12), .D(n46_adj_257), 
         .Z(n20)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut.init = 16'hfefc;
    LUT4 Select_4290_i7_2_lut (.A(databus_out[7]), .B(rw), .Z(n7)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4290_i7_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_353 (.A(read_value[7]), .B(n14_c), .C(n3), .D(n46), 
         .Z(n18_c)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_353.init = 16'hfefc;
    LUT4 i1_4_lut (.A(read_value_adj_308[7]), .B(read_value_adj_310[7]), 
         .C(n52), .D(n64), .Z(n12)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i3_4_lut_adj_354 (.A(read_value_adj_309[7]), .B(n66), .C(n52_adj_158), 
         .D(read_value_adj_311[7]), .Z(n14_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_354.init = 16'heca0;
    LUT4 i14_2_lut (.A(\select[7] ), .B(rw), .Z(n46_adj_257)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(214[19:32])
    defparam i14_2_lut.init = 16'h8888;
    LUT4 Select_4271_i5_2_lut (.A(databus_out[14]), .B(rw), .Z(n5_adj_263)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4271_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_355 (.A(read_value_adj_309[14]), .B(\read_value[14]_adj_190 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_265)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_355.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_22706 (.A(\register[6] [6]), .B(\register_addr[0] ), 
         .Z(n30816)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22706.init = 16'h2222;
    LUT4 i10_4_lut_adj_356 (.A(n15_adj_266), .B(n20_adj_267), .C(n2_adj_191), 
         .D(n7_adj_269), .Z(databus[6])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_356.init = 16'hfffe;
    LUT4 register_addr_1__bdd_3_lut_22707 (.A(\register_addr[0] ), .B(\register[4] [6]), 
         .C(\register[5] [6]), .Z(n30817)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22707.init = 16'he4e4;
    LUT4 i4_4_lut_adj_357 (.A(\read_value[6]_adj_192 ), .B(\read_value[6]_adj_193 ), 
         .C(n31447), .D(n31444), .Z(n15_adj_266)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_357.init = 16'heca0;
    LUT4 i9_4_lut_adj_358 (.A(read_value_adj_588[6]), .B(n18_adj_272), .C(n12_adj_273), 
         .D(n46_adj_257), .Z(n20_adj_267)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_358.init = 16'hfefc;
    LUT4 Select_4291_i7_2_lut (.A(databus_out[6]), .B(rw), .Z(n7_adj_269)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4291_i7_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_359 (.A(read_value[6]), .B(n14_adj_275), .C(n3_adj_194), 
         .D(n46), .Z(n18_adj_272)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_359.init = 16'hfefc;
    LUT4 i1_4_lut_adj_360 (.A(read_value_adj_308[6]), .B(read_value_adj_310[6]), 
         .C(n52), .D(n64), .Z(n12_adj_273)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_360.init = 16'heca0;
    LUT4 i3_4_lut_adj_361 (.A(read_value_adj_309[6]), .B(n66), .C(n52_adj_158), 
         .D(read_value_adj_311[6]), .Z(n14_adj_275)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_361.init = 16'heca0;
    LUT4 n1225_bdd_3_lut_22701 (.A(\register[2] [6]), .B(\register[3] [6]), 
         .C(\register_addr[0] ), .Z(n30819)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1225_bdd_3_lut_22701.init = 16'hcaca;
    LUT4 i10_4_lut_adj_362 (.A(n15_adj_281), .B(n20_adj_282), .C(n2_adj_195), 
         .D(n7_adj_284), .Z(databus[5])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_362.init = 16'hfffe;
    LUT4 i4_4_lut_adj_363 (.A(\read_value[5]_adj_196 ), .B(\read_value[5]_adj_197 ), 
         .C(n31447), .D(n31444), .Z(n15_adj_281)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_363.init = 16'heca0;
    LUT4 i9_4_lut_adj_364 (.A(read_value_adj_588[5]), .B(n18_adj_287), .C(n12_adj_288), 
         .D(n46_adj_257), .Z(n20_adj_282)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_364.init = 16'hfefc;
    LUT4 Select_4292_i7_2_lut (.A(databus_out[5]), .B(n33385), .Z(n7_adj_284)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4292_i7_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_365 (.A(read_value[5]), .B(n14_adj_290), .C(n3_adj_198), 
         .D(n46), .Z(n18_adj_287)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_365.init = 16'hfefc;
    LUT4 i1_4_lut_adj_366 (.A(read_value_adj_308[5]), .B(read_value_adj_310[5]), 
         .C(n52), .D(n64), .Z(n12_adj_288)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_366.init = 16'heca0;
    LUT4 i3_4_lut_adj_367 (.A(read_value_adj_309[5]), .B(n66), .C(n52_adj_158), 
         .D(read_value_adj_311[5]), .Z(n14_adj_290)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_367.init = 16'heca0;
    LUT4 n1225_bdd_3_lut_22964 (.A(n1225), .B(\register_addr[0] ), .C(\register[1] [6]), 
         .Z(n30820)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1225_bdd_3_lut_22964.init = 16'he2e2;
    LUT4 i10_4_lut_adj_368 (.A(n15_adj_296), .B(n20_adj_297), .C(n2_adj_199), 
         .D(n7_adj_299), .Z(databus[4])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_368.init = 16'hfffe;
    LUT4 i4_4_lut_adj_369 (.A(\read_value[4]_adj_200 ), .B(\read_value[4]_adj_201 ), 
         .C(n31447), .D(n31444), .Z(n15_adj_296)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_369.init = 16'heca0;
    LUT4 i9_4_lut_adj_370 (.A(read_value_adj_588[4]), .B(n18_adj_302), .C(n12_adj_303), 
         .D(n46_adj_257), .Z(n20_adj_297)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_370.init = 16'hfefc;
    LUT4 n1240_bdd_3_lut_22872 (.A(\register[2] [7]), .B(\register[3] [7]), 
         .C(\register_addr[0] ), .Z(n31157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1240_bdd_3_lut_22872.init = 16'hcaca;
    LUT4 Select_4293_i7_2_lut (.A(databus_out[4]), .B(n33385), .Z(n7_adj_299)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4293_i7_2_lut.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut_22930 (.A(\register_addr[0] ), .B(\register[4] [7]), 
         .C(\register[5] [7]), .Z(n31155)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22930.init = 16'he4e4;
    LUT4 n1240_bdd_3_lut_23346 (.A(n1240), .B(\register_addr[0] ), .C(\register[1] [7]), 
         .Z(n31158)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1240_bdd_3_lut_23346.init = 16'he2e2;
    LUT4 register_addr_1__bdd_2_lut_22929 (.A(\register[6] [7]), .B(\register_addr[0] ), 
         .Z(n31154)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22929.init = 16'h2222;
    LUT4 i7_4_lut_adj_371 (.A(read_value[4]), .B(n14_adj_305), .C(n3_adj_202), 
         .D(n46), .Z(n18_adj_302)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_371.init = 16'hfefc;
    LUT4 i1_4_lut_adj_372 (.A(read_value_adj_308[4]), .B(read_value_adj_310[4]), 
         .C(n52), .D(n64), .Z(n12_adj_303)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_372.init = 16'heca0;
    LUT4 i3_4_lut_adj_373 (.A(read_value_adj_309[4]), .B(read_value_adj_311[4]), 
         .C(n52_adj_158), .D(n66), .Z(n14_adj_305)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_373.init = 16'heca0;
    LUT4 i10_4_lut_adj_374 (.A(n15_adj_311), .B(n20_adj_312), .C(n2_adj_203), 
         .D(n7_adj_314), .Z(databus[3])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_374.init = 16'hfffe;
    LUT4 i4_4_lut_adj_375 (.A(\read_value[3]_adj_204 ), .B(\read_value[3]_adj_205 ), 
         .C(n31447), .D(n31444), .Z(n15_adj_311)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_375.init = 16'heca0;
    LUT4 i9_4_lut_adj_376 (.A(read_value_adj_588[3]), .B(n18_adj_317), .C(n12_adj_318), 
         .D(n46_adj_257), .Z(n20_adj_312)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_376.init = 16'hfefc;
    LUT4 i7_4_lut_adj_377 (.A(n13_adj_319), .B(n11_adj_320), .C(n2_adj_206), 
         .D(n5_adj_322), .Z(databus[22])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_377.init = 16'hfffe;
    LUT4 i5_4_lut_adj_378 (.A(\read_value[22]_adj_207 ), .B(n10_adj_323), 
         .C(n8_adj_208), .D(n31426), .Z(n13_adj_319)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_378.init = 16'hfefc;
    LUT4 i3_4_lut_adj_379 (.A(read_value[22]), .B(read_value_adj_308[22]), 
         .C(n46), .D(n52), .Z(n11_adj_320)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_379.init = 16'heca0;
    LUT4 Select_4294_i7_2_lut (.A(databus_out[3]), .B(n33385), .Z(n7_adj_314)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4294_i7_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_380 (.A(read_value[3]), .B(n14_adj_328), .C(n3_adj_209), 
         .D(n46), .Z(n18_adj_317)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_380.init = 16'hfefc;
    LUT4 i1_4_lut_adj_381 (.A(read_value_adj_308[3]), .B(read_value_adj_310[3]), 
         .C(n52), .D(n64), .Z(n12_adj_318)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_381.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_22743 (.A(\register[6] [2]), .B(\register_addr[0] ), 
         .Z(n30838)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22743.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut_22744 (.A(\register_addr[0] ), .B(\register[4] [2]), 
         .C(\register[5] [2]), .Z(n30839)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22744.init = 16'he4e4;
    LUT4 i3_4_lut_adj_382 (.A(read_value_adj_309[3]), .B(read_value_adj_311[3]), 
         .C(n52_adj_158), .D(n66), .Z(n14_adj_328)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_382.init = 16'heca0;
    LUT4 i10_4_lut_adj_383 (.A(n15_adj_334), .B(n20_adj_335), .C(n2_adj_210), 
         .D(n7_adj_337), .Z(databus[2])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_383.init = 16'hfffe;
    LUT4 n1195_bdd_3_lut_22716 (.A(\register[2] [2]), .B(\register[3] [2]), 
         .C(\register_addr[0] ), .Z(n30841)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1195_bdd_3_lut_22716.init = 16'hcaca;
    LUT4 Select_4247_i5_2_lut (.A(databus_out[22]), .B(rw), .Z(n5_adj_322)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4247_i5_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_384 (.A(\read_value[2]_adj_211 ), .B(\read_value[2]_adj_212 ), 
         .C(n31447), .D(n31444), .Z(n15_adj_334)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_384.init = 16'heca0;
    LUT4 i9_4_lut_adj_385 (.A(read_value_adj_588[2]), .B(n18_adj_340), .C(n12_adj_341), 
         .D(n46_adj_257), .Z(n20_adj_335)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_385.init = 16'hfefc;
    LUT4 Select_4295_i7_2_lut (.A(databus_out[2]), .B(n33385), .Z(n7_adj_337)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4295_i7_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_386 (.A(read_value_adj_309[22]), .B(\read_value[22]_adj_213 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_323)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_386.init = 16'heca0;
    LUT4 i7_4_lut_adj_387 (.A(read_value[2]), .B(n14_adj_345), .C(n3_adj_214), 
         .D(n46), .Z(n18_adj_340)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_387.init = 16'hfefc;
    LUT4 i1_4_lut_adj_388 (.A(read_value_adj_308[2]), .B(read_value_adj_310[2]), 
         .C(n52), .D(n64), .Z(n12_adj_341)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_388.init = 16'heca0;
    LUT4 i3_4_lut_adj_389 (.A(read_value_adj_309[2]), .B(read_value_adj_311[2]), 
         .C(n52_adj_158), .D(n66), .Z(n14_adj_345)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_389.init = 16'heca0;
    LUT4 n1195_bdd_3_lut_22941 (.A(n1195), .B(\register_addr[0] ), .C(\register[1] [2]), 
         .Z(n30842)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1195_bdd_3_lut_22941.init = 16'he2e2;
    LUT4 i10_4_lut_adj_390 (.A(n19), .B(n8_adj_351), .C(n18_adj_352), 
         .D(n12_adj_353), .Z(databus[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_390.init = 16'hfffe;
    LUT4 i8_4_lut (.A(read_value_adj_588[1]), .B(n16), .C(n10), .D(n46_adj_257), 
         .Z(n19)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut.init = 16'hfefc;
    LUT4 Select_4296_i8_2_lut (.A(databus_out[1]), .B(rw), .Z(n8_adj_351)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4296_i8_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_391 (.A(\read_value[1]_adj_215 ), .B(n14_adj_356), 
         .C(n3_adj_216), .D(n31444), .Z(n18_adj_352)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_391.init = 16'hfefc;
    LUT4 i1_4_lut_adj_392 (.A(read_value_adj_308[1]), .B(read_value_adj_310[1]), 
         .C(n52), .D(n64), .Z(n12_adj_353)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_392.init = 16'heca0;
    LUT4 i5_4_lut_adj_393 (.A(\read_value[1]_adj_217 ), .B(read_value[1]), 
         .C(n31426), .D(n46), .Z(n16)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i5_4_lut_adj_393.init = 16'heca0;
    LUT4 i3_4_lut_adj_394 (.A(read_value_adj_309[1]), .B(read_value_adj_311[1]), 
         .C(n52_adj_158), .D(n66), .Z(n14_adj_356)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_394.init = 16'heca0;
    LUT4 i7_4_lut_adj_395 (.A(n13_adj_364), .B(n11_adj_365), .C(n2_adj_218), 
         .D(n5_adj_367), .Z(databus[13])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_395.init = 16'hfffe;
    LUT4 i5_4_lut_adj_396 (.A(\read_value[13]_adj_219 ), .B(n10_adj_368), 
         .C(n8_adj_220), .D(n31426), .Z(n13_adj_364)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_396.init = 16'hfefc;
    LUT4 i7_4_lut_adj_397 (.A(n13_adj_370), .B(n11_adj_371), .C(n2_adj_221), 
         .D(n5_adj_373), .Z(databus[23])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_397.init = 16'hfffe;
    LUT4 i3_4_lut_adj_398 (.A(read_value[13]), .B(read_value_adj_308[13]), 
         .C(n46), .D(n52), .Z(n11_adj_365)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_398.init = 16'heca0;
    LUT4 Select_4274_i5_2_lut (.A(databus_out[13]), .B(n33385), .Z(n5_adj_367)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4274_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_399 (.A(read_value_adj_309[13]), .B(\read_value[13]_adj_222 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_368)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_399.init = 16'heca0;
    LUT4 i5_4_lut_adj_400 (.A(\read_value[23]_adj_223 ), .B(n10_adj_378), 
         .C(n8_adj_224), .D(n31426), .Z(n13_adj_370)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_400.init = 16'hfefc;
    LUT4 i3_4_lut_adj_401 (.A(read_value[23]), .B(read_value_adj_308[23]), 
         .C(n46), .D(n52), .Z(n11_adj_371)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_401.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_22585 (.A(\register_addr[0] ), .B(\register[4] [5]), 
         .C(\register[5] [5]), .Z(n30334)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22585.init = 16'he4e4;
    LUT4 i7_4_lut_adj_402 (.A(n13_adj_382), .B(n11_adj_383), .C(n2_adj_225), 
         .D(n5_adj_385), .Z(databus[21])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_402.init = 16'hfffe;
    LUT4 Select_4244_i5_2_lut (.A(databus_out[23]), .B(rw), .Z(n5_adj_373)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4244_i5_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_403 (.A(n13_adj_386), .B(n11_adj_387), .C(n2_adj_226), 
         .D(n5_adj_389), .Z(databus[12])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_403.init = 16'hfffe;
    LUT4 i5_4_lut_adj_404 (.A(\read_value[12]_adj_227 ), .B(n10_adj_390), 
         .C(n8_adj_228), .D(n31426), .Z(n13_adj_386)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_404.init = 16'hfefc;
    LUT4 i2_4_lut_adj_405 (.A(read_value_adj_309[23]), .B(\read_value[23]_adj_229 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_378)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_405.init = 16'heca0;
    LUT4 i3_4_lut_adj_406 (.A(read_value[12]), .B(read_value_adj_308[12]), 
         .C(n46), .D(n52), .Z(n11_adj_387)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_406.init = 16'heca0;
    LUT4 Select_4277_i5_2_lut (.A(databus_out[12]), .B(n33385), .Z(n5_adj_389)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4277_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_407 (.A(read_value_adj_309[12]), .B(\read_value[12]_adj_230 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_390)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_407.init = 16'heca0;
    LUT4 i5_4_lut_adj_408 (.A(\read_value[21]_adj_231 ), .B(n10_adj_398), 
         .C(n8_adj_232), .D(n31426), .Z(n13_adj_382)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_408.init = 16'hfefc;
    LUT4 i3_4_lut_adj_409 (.A(read_size[0]), .B(read_size_c[0]), .C(\select[1] ), 
         .D(\select[7] ), .Z(n13)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_409.init = 16'heca0;
    LUT4 i8_4_lut_adj_410 (.A(n31483), .B(n16_adj_402), .C(n9), .D(\read_size[0]_adj_233 ), 
         .Z(n18)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_410.init = 16'hfefc;
    LUT4 i4_4_lut_adj_411 (.A(\read_size[0]_adj_234 ), .B(\read_size[0]_adj_235 ), 
         .C(n31465), .D(\select[2] ), .Z(n14)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_411.init = 16'heca0;
    LUT4 i6_4_lut (.A(n31474), .B(n12_adj_408), .C(n5), .D(\read_size[0]_adj_236 ), 
         .Z(n16_adj_402)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut.init = 16'hfefc;
    LUT4 i3_4_lut_adj_412 (.A(read_value[21]), .B(read_value_adj_308[21]), 
         .C(n46), .D(n52), .Z(n11_adj_383)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_412.init = 16'heca0;
    LUT4 i2_4_lut_adj_413 (.A(\read_size[0]_adj_237 ), .B(n31445), .C(\select[5] ), 
         .D(\read_size[0]_adj_238 ), .Z(n12_adj_408)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_413.init = 16'heca0;
    LUT4 i7_4_lut_adj_414 (.A(n13_adj_415), .B(n11_adj_416), .C(n2_adj_239), 
         .D(n5_adj_418), .Z(databus[11])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_414.init = 16'hfffe;
    LUT4 i5_4_lut_adj_415 (.A(\read_value[11]_adj_240 ), .B(n10_adj_419), 
         .C(n8_adj_241), .D(n31426), .Z(n13_adj_415)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_415.init = 16'hfefc;
    LUT4 i3_4_lut_adj_416 (.A(read_value[11]), .B(read_value_adj_308[11]), 
         .C(n46), .D(n52), .Z(n11_adj_416)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_416.init = 16'heca0;
    LUT4 i5_4_lut_adj_417 (.A(n31445), .B(n10_adj_423), .C(n6), .D(\read_size[2]_adj_242 ), 
         .Z(\reg_size[2] )) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_417.init = 16'hfefc;
    LUT4 i4_4_lut_adj_418 (.A(\read_size[2]_adj_243 ), .B(n8_adj_425), .C(n9_adj_244), 
         .D(n31483), .Z(n10_adj_423)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_418.init = 16'hfefc;
    LUT4 n1180_bdd_3_lut_22749 (.A(\register[2] [1]), .B(\register[3] [1]), 
         .C(\register_addr[0] ), .Z(n30888)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1180_bdd_3_lut_22749.init = 16'hcaca;
    LUT4 i2_4_lut_adj_419 (.A(read_size[2]), .B(\read_size[2]_adj_245 ), 
         .C(\select[1] ), .D(n31471), .Z(n8_adj_425)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_419.init = 16'heca0;
    LUT4 Select_4280_i5_2_lut (.A(databus_out[11]), .B(n33385), .Z(n5_adj_418)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4280_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_420 (.A(read_value_adj_309[11]), .B(\read_value[11]_adj_246 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_419)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_420.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_22788 (.A(\register[6] [1]), .B(\register_addr[0] ), 
         .Z(n30885)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22788.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut_22789 (.A(\register_addr[0] ), .B(\register[4] [1]), 
         .C(\register[5] [1]), .Z(n30886)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22789.init = 16'he4e4;
    LUT4 n1180_bdd_3_lut_22913 (.A(n1180), .B(\register_addr[0] ), .C(\register[1] [1]), 
         .Z(n30889)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1180_bdd_3_lut_22913.init = 16'he2e2;
    LUT4 Select_4250_i5_2_lut (.A(databus_out[21]), .B(rw), .Z(n5_adj_385)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4250_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_421 (.A(read_value_adj_309[21]), .B(\read_value[21]_adj_247 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_398)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_421.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_22952 (.A(\register_addr[0] ), .B(\register[4] [4]), 
         .C(\register[5] [4]), .Z(n31305)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_22952.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_22951 (.A(\register[6] [4]), .B(\register_addr[0] ), 
         .Z(n31304)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_22951.init = 16'h2222;
    LUT4 \register_1[[4__bdd_3_lut_23198  (.A(\register[2] [4]), .B(\register[3] [4]), 
         .C(\register_addr[0] ), .Z(n31307)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[4__bdd_3_lut_23198 .init = 16'hcaca;
    LUT4 \register_1[[4__bdd_2_lut_23199  (.A(\register[1] [4]), .B(\register_addr[0] ), 
         .Z(n31308)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[4__bdd_2_lut_23199 .init = 16'h8888;
    LUT4 i7_4_lut_adj_422 (.A(n13_adj_433), .B(n11_adj_434), .C(n2_adj_248), 
         .D(n5_adj_436), .Z(databus[25])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_422.init = 16'hfffe;
    LUT4 register_addr_1__bdd_3_lut (.A(\register_addr[0] ), .B(\register[4] [0]), 
         .C(\register[5] [0]), .Z(n31317)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut.init = 16'he4e4;
    LUT4 i5_4_lut_adj_423 (.A(\read_value[25]_adj_249 ), .B(n10_adj_437), 
         .C(n8_adj_250), .D(n31426), .Z(n13_adj_433)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_423.init = 16'hfefc;
    LUT4 i3_4_lut_adj_424 (.A(read_value[25]), .B(read_value_adj_308[25]), 
         .C(n46), .D(n52), .Z(n11_adj_434)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_424.init = 16'heca0;
    LUT4 Select_4238_i5_2_lut (.A(databus_out[25]), .B(rw), .Z(n5_adj_436)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4238_i5_2_lut.init = 16'h2222;
    LUT4 register_addr_1__bdd_2_lut (.A(\register[6] [0]), .B(\register_addr[0] ), 
         .Z(n31316)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_425 (.A(read_value_adj_309[25]), .B(\read_value[25]_adj_251 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_437)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_425.init = 16'heca0;
    L6MUX21 i22958 (.D0(n31321), .D1(n31318), .SD(\register_addr[2] ), 
            .Z(n31322));
    LUT4 n1165_bdd_3_lut_22955 (.A(\register[2] [0]), .B(\register[3] [0]), 
         .C(\register_addr[0] ), .Z(n31319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1165_bdd_3_lut_22955.init = 16'hcaca;
    PFUMX i22956 (.BLUT(n31320), .ALUT(n31319), .C0(\register_addr[1] ), 
          .Z(n31321));
    LUT4 n1165_bdd_3_lut_23162 (.A(n1165), .B(\register_addr[0] ), .C(\register[1] [0]), 
         .Z(n31320)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1165_bdd_3_lut_23162.init = 16'he2e2;
    LUT4 i7_4_lut_adj_426 (.A(n13_adj_443), .B(n11_adj_444), .C(n2_adj_252), 
         .D(n5_adj_446), .Z(databus[20])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_426.init = 16'hfffe;
    PFUMX i22953 (.BLUT(n31317), .ALUT(n31316), .C0(\register_addr[1] ), 
          .Z(n31318));
    LUT4 i7_4_lut_adj_427 (.A(n13_adj_447), .B(n11_adj_448), .C(n2_adj_253), 
         .D(n5_adj_450), .Z(databus[16])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_427.init = 16'hfffe;
    LUT4 i5_4_lut_adj_428 (.A(\read_value[20]_adj_254 ), .B(n10_adj_451), 
         .C(n8_adj_255), .D(n31426), .Z(n13_adj_443)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_428.init = 16'hfefc;
    LUT4 i5_4_lut_adj_429 (.A(\read_value[16]_adj_256 ), .B(n10_adj_453), 
         .C(n8_adj_257), .D(n31426), .Z(n13_adj_447)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_429.init = 16'hfefc;
    L6MUX21 i22949 (.D0(n31309), .D1(n31306), .SD(\register_addr[2] ), 
            .Z(n31310));
    PFUMX i22947 (.BLUT(n31308), .ALUT(n31307), .C0(\register_addr[1] ), 
          .Z(n31309));
    LUT4 i3_4_lut_adj_430 (.A(read_value[20]), .B(read_value_adj_308[20]), 
         .C(n46), .D(n52), .Z(n11_adj_444)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_430.init = 16'heca0;
    LUT4 Select_4307_i1_2_lut_rep_444 (.A(read_size[1]), .B(\select[1] ), 
         .Z(n31588)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4307_i1_2_lut_rep_444.init = 16'h8888;
    LUT4 i3_4_lut_adj_431 (.A(read_value[16]), .B(read_value_adj_308[16]), 
         .C(n46), .D(n52), .Z(n11_adj_448)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_431.init = 16'heca0;
    LUT4 i1_2_lut_3_lut (.A(read_size[1]), .B(\select[1] ), .C(\sendcount[1] ), 
         .Z(n13156)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7878;
    LUT4 Select_4265_i5_2_lut (.A(databus_out[16]), .B(n33385), .Z(n5_adj_450)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4265_i5_2_lut.init = 16'h2222;
    FD1S3IX read_value__i1 (.D(n30891), .CK(\select[7] ), .CD(n31457), 
            .Q(read_value_adj_588[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1S3IX read_value__i2 (.D(n30844), .CK(\select[7] ), .CD(n31457), 
            .Q(read_value_adj_588[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1S3IX read_value__i3 (.D(n30783), .CK(\select[7] ), .CD(n31457), 
            .Q(read_value_adj_588[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1S3IX read_value__i4 (.D(n31310), .CK(\select[7] ), .CD(n31457), 
            .Q(read_value_adj_588[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1S3IX read_value__i5 (.D(n30339), .CK(\select[7] ), .CD(n31457), 
            .Q(read_value_adj_588[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1S3IX read_value__i6 (.D(n30822), .CK(\select[7] ), .CD(n31457), 
            .Q(read_value_adj_588[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1S3IX read_value__i7 (.D(n31160), .CK(\select[7] ), .CD(n31457), 
            .Q(read_value_adj_588[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i7.GSR = "ENABLED";
    PFUMX i22945 (.BLUT(n31305), .ALUT(n31304), .C0(\register_addr[1] ), 
          .Z(n31306));
    LUT4 Select_4253_i5_2_lut (.A(databus_out[20]), .B(rw), .Z(n5_adj_446)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4253_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_432 (.A(read_value_adj_309[20]), .B(\read_value[20]_adj_258 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_451)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_432.init = 16'heca0;
    LUT4 i7_4_lut_adj_433 (.A(n13_adj_461), .B(n11_adj_462), .C(n2_adj_259), 
         .D(n5_adj_263), .Z(databus[14])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_433.init = 16'hfffe;
    LUT4 i10_4_lut_adj_434 (.A(n15_adj_464), .B(n20_adj_465), .C(n2_adj_260), 
         .D(n7_adj_467), .Z(databus[0])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_434.init = 16'hfffe;
    LUT4 i4_4_lut_adj_435 (.A(\read_value[0]_adj_261 ), .B(\read_value[0]_adj_262 ), 
         .C(n31447), .D(n31444), .Z(n15_adj_464)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_435.init = 16'heca0;
    LUT4 i9_4_lut_adj_436 (.A(read_value_adj_588[0]), .B(n18_adj_470), .C(n12_adj_471), 
         .D(n46_adj_257), .Z(n20_adj_465)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_436.init = 16'hfefc;
    LUT4 Select_4297_i7_2_lut (.A(databus_out[0]), .B(rw), .Z(n7_adj_467)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4297_i7_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_437 (.A(read_value[0]), .B(n14_adj_473), .C(n3_adj_263), 
         .D(n46), .Z(n18_adj_470)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_437.init = 16'hfefc;
    LUT4 i7_4_lut_adj_438 (.A(n13_adj_475), .B(n11_adj_476), .C(n2_adj_264), 
         .D(n5_adj_478), .Z(databus[26])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_438.init = 16'hfffe;
    LUT4 i1_4_lut_adj_439 (.A(read_value_adj_308[0]), .B(read_value_adj_310[0]), 
         .C(n52), .D(n64), .Z(n12_adj_471)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_439.init = 16'heca0;
    LUT4 i5_4_lut_adj_440 (.A(\read_value[26]_adj_265 ), .B(n10_adj_481), 
         .C(n8_adj_266), .D(n31426), .Z(n13_adj_475)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_440.init = 16'hfefc;
    LUT4 i3_4_lut_adj_441 (.A(read_value_adj_309[0]), .B(n66), .C(n52_adj_158), 
         .D(read_value_adj_311[0]), .Z(n14_adj_473)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_441.init = 16'heca0;
    LUT4 i3_4_lut_adj_442 (.A(read_value[26]), .B(read_value_adj_308[26]), 
         .C(n46), .D(n52), .Z(n11_adj_476)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_442.init = 16'heca0;
    LUT4 Select_4235_i5_2_lut (.A(databus_out[26]), .B(rw), .Z(n5_adj_478)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4235_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_443 (.A(read_value_adj_309[26]), .B(\read_value[26]_adj_267 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_481)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_443.init = 16'heca0;
    LUT4 i2_4_lut_adj_444 (.A(read_value_adj_309[16]), .B(\read_value[16]_adj_268 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_453)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_444.init = 16'heca0;
    L6MUX21 i22583 (.D0(n30338), .D1(n30335), .SD(\register_addr[2] ), 
            .Z(n30339));
    L6MUX21 i22875 (.D0(n31159), .D1(n31156), .SD(\register_addr[2] ), 
            .Z(n31160));
    PFUMX i22873 (.BLUT(n31158), .ALUT(n31157), .C0(\register_addr[1] ), 
          .Z(n31159));
    LUT4 i7_4_lut_adj_445 (.A(n13_adj_491), .B(n11_adj_492), .C(n2_adj_269), 
         .D(n5_adj_494), .Z(databus[19])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_445.init = 16'hfffe;
    PFUMX i22870 (.BLUT(n31155), .ALUT(n31154), .C0(\register_addr[1] ), 
          .Z(n31156));
    LUT4 i5_4_lut_adj_446 (.A(\read_value[19]_adj_270 ), .B(n10_adj_495), 
         .C(n8_adj_271), .D(n31426), .Z(n13_adj_491)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_446.init = 16'hfefc;
    LUT4 i1_2_lut (.A(\register_addr[0] ), .B(\register_addr[1] ), .Z(n29237)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    PFUMX i22581 (.BLUT(n30337), .ALUT(n30336), .C0(\register_addr[1] ), 
          .Z(n30338));
    LUT4 i3_4_lut_adj_447 (.A(read_value[19]), .B(read_value_adj_308[19]), 
         .C(n46), .D(n52), .Z(n11_adj_492)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_447.init = 16'heca0;
    FD1S3IX read_value__i0 (.D(n31322), .CK(\select[7] ), .CD(n31457), 
            .Q(read_value_adj_588[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i7_4_lut_adj_448 (.A(n13_adj_499), .B(n11_adj_500), .C(n2_adj_272), 
         .D(n5_adj_502), .Z(databus[15])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_448.init = 16'hfffe;
    LUT4 Select_4256_i5_2_lut (.A(databus_out[19]), .B(rw), .Z(n5_adj_494)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4256_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_449 (.A(read_value_adj_309[19]), .B(\read_value[19]_adj_273 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_495)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_449.init = 16'heca0;
    L6MUX21 i22752 (.D0(n30890), .D1(n30887), .SD(\register_addr[2] ), 
            .Z(n30891));
    PFUMX i22750 (.BLUT(n30889), .ALUT(n30888), .C0(\register_addr[1] ), 
          .Z(n30890));
    LUT4 i7_4_lut_adj_450 (.A(n13_adj_505), .B(n11_adj_506), .C(n2_adj_274), 
         .D(n5_adj_508), .Z(databus[18])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_450.init = 16'hfffe;
    LUT4 i5_4_lut_adj_451 (.A(\read_value[18]_adj_275 ), .B(n10_adj_509), 
         .C(n8_adj_276), .D(n31426), .Z(n13_adj_505)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_451.init = 16'hfefc;
    LUT4 i3_4_lut_adj_452 (.A(read_value[18]), .B(read_value_adj_308[18]), 
         .C(n46), .D(n52), .Z(n11_adj_506)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_452.init = 16'heca0;
    PFUMX i22747 (.BLUT(n30886), .ALUT(n30885), .C0(\register_addr[1] ), 
          .Z(n30887));
    LUT4 i7_4_lut_adj_453 (.A(n13_adj_513), .B(n11_adj_514), .C(n2_adj_277), 
         .D(n5_adj_516), .Z(databus[31])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_453.init = 16'hfffe;
    LUT4 i5_4_lut_adj_454 (.A(\read_value[31]_adj_278 ), .B(n10_adj_517), 
         .C(n8_adj_279), .D(n31426), .Z(n13_adj_513)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_454.init = 16'hfefc;
    LUT4 i3_4_lut_adj_455 (.A(read_value[31]), .B(read_value_adj_308[31]), 
         .C(n46), .D(n52), .Z(n11_adj_514)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_455.init = 16'heca0;
    LUT4 Select_4262_i5_2_lut (.A(databus_out[17]), .B(n33385), .Z(n5_adj_521)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4262_i5_2_lut.init = 16'h2222;
    LUT4 i5_4_lut_adj_456 (.A(\read_value[14]_adj_280 ), .B(n10_adj_265), 
         .C(n8_adj_281), .D(n31426), .Z(n13_adj_461)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_456.init = 16'hfefc;
    LUT4 Select_4259_i5_2_lut (.A(databus_out[18]), .B(n33385), .Z(n5_adj_508)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4259_i5_2_lut.init = 16'h2222;
    LUT4 Select_4220_i5_2_lut (.A(databus_out[31]), .B(rw), .Z(n5_adj_516)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4220_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_457 (.A(read_value_adj_309[31]), .B(\read_value[31]_adj_282 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_517)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_457.init = 16'heca0;
    LUT4 i7_4_lut_adj_458 (.A(n13_adj_526), .B(n11_adj_527), .C(n2_adj_283), 
         .D(n5_adj_529), .Z(databus[30])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_458.init = 16'hfffe;
    LUT4 i5_4_lut_adj_459 (.A(\read_value[30]_adj_284 ), .B(n10_adj_530), 
         .C(n8_adj_285), .D(n31426), .Z(n13_adj_526)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_459.init = 16'hfefc;
    L6MUX21 i22719 (.D0(n30843), .D1(n30840), .SD(\register_addr[2] ), 
            .Z(n30844));
    LUT4 i3_4_lut_adj_460 (.A(read_value[30]), .B(read_value_adj_308[30]), 
         .C(n46), .D(n52), .Z(n11_adj_527)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_460.init = 16'heca0;
    LUT4 i2_4_lut_adj_461 (.A(read_value_adj_309[18]), .B(\read_value[18]_adj_286 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_509)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_461.init = 16'heca0;
    LUT4 Select_4223_i5_2_lut (.A(databus_out[30]), .B(rw), .Z(n5_adj_529)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4223_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_462 (.A(read_value_adj_309[30]), .B(\read_value[30]_adj_287 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_530)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_462.init = 16'heca0;
    PFUMX i22717 (.BLUT(n30842), .ALUT(n30841), .C0(\register_addr[1] ), 
          .Z(n30843));
    LUT4 \register_1[[5__bdd_3_lut_22781  (.A(\register[2] [5]), .B(\register[3] [5]), 
         .C(\register_addr[0] ), .Z(n30336)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[5__bdd_3_lut_22781 .init = 16'hcaca;
    LUT4 i7_4_lut_adj_463 (.A(n13_adj_538), .B(n11_adj_539), .C(n2_adj_288), 
         .D(n5_adj_541), .Z(databus[29])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_463.init = 16'hfffe;
    LUT4 i2_4_lut_adj_464 (.A(read_value_adj_309[17]), .B(\read_value[17]_adj_289 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_543)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_464.init = 16'heca0;
    LUT4 i5_4_lut_adj_465 (.A(\read_value[29]_adj_290 ), .B(n10_adj_544), 
         .C(n8_adj_291), .D(n31426), .Z(n13_adj_538)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_465.init = 16'hfefc;
    LUT4 i3_4_lut_adj_466 (.A(read_value[29]), .B(read_value_adj_308[29]), 
         .C(n46), .D(n52), .Z(n11_adj_539)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_466.init = 16'heca0;
    LUT4 Select_4226_i5_2_lut (.A(databus_out[29]), .B(rw), .Z(n5_adj_541)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4226_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_467 (.A(read_value_adj_309[29]), .B(\read_value[29]_adj_292 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_544)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_467.init = 16'heca0;
    PFUMX i22714 (.BLUT(n30839), .ALUT(n30838), .C0(\register_addr[1] ), 
          .Z(n30840));
    LUT4 i7_4_lut_adj_468 (.A(n13_adj_550), .B(n11_adj_551), .C(n2_adj_293), 
         .D(n5_adj_553), .Z(databus[28])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_468.init = 16'hfffe;
    LUT4 i3_4_lut_adj_469 (.A(read_value[14]), .B(read_value_adj_308[14]), 
         .C(n46), .D(n52), .Z(n11_adj_462)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_469.init = 16'heca0;
    LUT4 i7_4_lut_adj_470 (.A(n13_adj_556), .B(n11_adj_557), .C(n2_adj_294), 
         .D(n5_adj_521), .Z(databus[17])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_470.init = 16'hfffe;
    LUT4 i5_4_lut_adj_471 (.A(\read_value[15]_adj_295 ), .B(n10_adj_559), 
         .C(n8_adj_296), .D(n31426), .Z(n13_adj_499)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_471.init = 16'hfefc;
    L6MUX21 i22704 (.D0(n30821), .D1(n30818), .SD(\register_addr[2] ), 
            .Z(n30822));
    LUT4 i3_4_lut_adj_472 (.A(read_value[15]), .B(read_value_adj_308[15]), 
         .C(n46), .D(n52), .Z(n11_adj_500)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_472.init = 16'heca0;
    PFUMX i22702 (.BLUT(n30820), .ALUT(n30819), .C0(\register_addr[1] ), 
          .Z(n30821));
    PFUMX i22699 (.BLUT(n30817), .ALUT(n30816), .C0(\register_addr[1] ), 
          .Z(n30818));
    LUT4 i5_4_lut_adj_473 (.A(\read_value[28]_adj_297 ), .B(n10_adj_563), 
         .C(n8_adj_298), .D(n31426), .Z(n13_adj_550)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_473.init = 16'hfefc;
    LUT4 i3_4_lut_adj_474 (.A(read_value[28]), .B(read_value_adj_308[28]), 
         .C(n46), .D(n52), .Z(n11_adj_551)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_474.init = 16'heca0;
    LUT4 Select_4229_i5_2_lut (.A(databus_out[28]), .B(rw), .Z(n5_adj_553)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4229_i5_2_lut.init = 16'h2222;
    LUT4 i5_4_lut_adj_475 (.A(\read_value[17]_adj_299 ), .B(n10_adj_543), 
         .C(n8_adj_300), .D(n31426), .Z(n13_adj_556)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_475.init = 16'hfefc;
    LUT4 i2_4_lut_adj_476 (.A(read_value_adj_309[28]), .B(\read_value[28]_adj_301 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_563)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_476.init = 16'heca0;
    PFUMX i22579 (.BLUT(n30334), .ALUT(n30333), .C0(\register_addr[1] ), 
          .Z(n30335));
    LUT4 i7_4_lut_adj_477 (.A(n13_adj_571), .B(n11_adj_572), .C(n2_adj_302), 
         .D(n5_adj_574), .Z(databus[27])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_477.init = 16'hfffe;
    LUT4 i5_4_lut_adj_478 (.A(\read_value[27]_adj_303 ), .B(n10_adj_575), 
         .C(n8_adj_304), .D(n31426), .Z(n13_adj_571)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_478.init = 16'hfefc;
    LUT4 i3_4_lut_adj_479 (.A(read_value[27]), .B(read_value_adj_308[27]), 
         .C(n46), .D(n52), .Z(n11_adj_572)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_479.init = 16'heca0;
    L6MUX21 i22683 (.D0(n30782), .D1(n30779), .SD(\register_addr[2] ), 
            .Z(n30783));
    LUT4 i3_4_lut_adj_480 (.A(read_value[17]), .B(read_value_adj_308[17]), 
         .C(n46), .D(n52), .Z(n11_adj_557)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_480.init = 16'heca0;
    LUT4 Select_4268_i5_2_lut (.A(databus_out[15]), .B(n33385), .Z(n5_adj_502)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4268_i5_2_lut.init = 16'h2222;
    PFUMX i22681 (.BLUT(n30781), .ALUT(n30780), .C0(\register_addr[1] ), 
          .Z(n30782));
    LUT4 Select_4232_i5_2_lut (.A(databus_out[27]), .B(rw), .Z(n5_adj_574)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4232_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_481 (.A(read_value_adj_309[15]), .B(\read_value[15]_adj_305 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_559)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_481.init = 16'heca0;
    LUT4 i2_4_lut_adj_482 (.A(read_value_adj_309[27]), .B(\read_value[27]_adj_306 ), 
         .C(n52_adj_158), .D(n31447), .Z(n10_adj_575)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_482.init = 16'heca0;
    PWMReceiver recv_ch8 (.GND_net(GND_net), .debug_c_c(debug_c_c), .n33387(n33387), 
            .rc_ch8_c(rc_ch8_c), .n29818(n29818), .n33386(n33386), .\register[6] ({\register[6] }), 
            .n13957(n13957), .n1240(n1240), .n27564(n27564), .n29784(n29784)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(257[14] 261[36])
    PWMReceiver_U1 recv_ch7 (.\register[5] ({\register[5] }), .debug_c_c(debug_c_c), 
            .n33386(n33386), .n33387(n33387), .rc_ch7_c(rc_ch7_c), .GND_net(GND_net), 
            .n33388(n33388), .n1225(n1225), .n27543(n27543), .n29827(n29827)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(252[14] 256[36])
    PWMReceiver_U2 recv_ch4 (.n33386(n33386), .debug_c_c(debug_c_c), .n33387(n33387), 
            .rc_ch4_c(rc_ch4_c), .GND_net(GND_net), .n33388(n33388), .\register[4] ({\register[4] }), 
            .n1210(n1210), .n27550(n27550), .n29838(n29838)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(247[14] 251[36])
    PWMReceiver_U3 recv_ch3 (.debug_c_c(debug_c_c), .n33387(n33387), .rc_ch3_c(rc_ch3_c), 
            .GND_net(GND_net), .n33388(n33388), .\register[3] ({\register[3] }), 
            .n14500(n14500), .n1195(n1195), .n27541(n27541), .n29840(n29840), 
            .n29530(n29530), .n29944(n29944), .n14(n14_adj_307)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(242[14] 246[36])
    PWMReceiver_U4 recv_ch2 (.GND_net(GND_net), .n29832(n29832), .debug_c_c(debug_c_c), 
            .n33387(n33387), .rc_ch2_c(rc_ch2_c), .n31412(n31412), .n33388(n33388), 
            .\register[2] ({\register[2] }), .n14513(n14513), .n29847(n29847), 
            .n1180(n1180), .n27536(n27536), .n33386(n33386), .n31512(n31512)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(237[14] 241[36])
    PWMReceiver_U5 recv_ch1 (.debug_c_c(debug_c_c), .n33387(n33387), .\register[1] ({\register[1] }), 
            .n14514(n14514), .rc_ch1_c(rc_ch1_c), .GND_net(GND_net), .n29830(n29830), 
            .n33386(n33386), .n1165(n1165), .n27547(n27547), .n29811(n29811)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(232[17] 236[36])
    
endmodule
//
// Verilog Description of module PWMReceiver
//

module PWMReceiver (GND_net, debug_c_c, n33387, rc_ch8_c, n29818, 
            n33386, \register[6] , n13957, n1240, n27564, n29784) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    input n33387;
    input rc_ch8_c;
    output n29818;
    input n33386;
    output [7:0]\register[6] ;
    input n13957;
    output n1240;
    input n27564;
    output n29784;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n27592, n31467, n31594, n31531, n27756, n31500, n27724, 
        n27395, n10, n26460, n31602;
    wire [15:0]n116;
    
    wire n26461, n31593, n29377, n31480, n1246, n1234, n31543, 
        n26459, n29253, n4, n26458, n26457, n31468, n26456, n29400, 
        n29314, n54, n29554, n23, n28997, n17066, n24;
    wire [7:0]n1138;
    wire [7:0]n43;
    
    wire n31597, n29472, n31532, n29250, n31583, n6, n31595, n4_adj_218, 
        n29401, n26463, n26462, n28988, n29562, n29638, n26735, 
        n26734, n26733, n26732;
    
    LUT4 i15626_2_lut_rep_323 (.A(count[9]), .B(n27592), .Z(n31467)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i15626_2_lut_rep_323.init = 16'h8888;
    LUT4 i2_3_lut_4_lut (.A(count[9]), .B(n27592), .C(n31594), .D(n31531), 
         .Z(n27756)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_3_lut_4_lut.init = 16'hfff8;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n31500), .C(n27724), 
         .D(n27395), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    CCU2D add_1795_11 (.A0(count[9]), .B0(n31602), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n31602), .C1(GND_net), .D1(GND_net), .CIN(n26460), 
          .COUT(n26461), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1795_11.INIT0 = 16'hd222;
    defparam add_1795_11.INIT1 = 16'hd222;
    defparam add_1795_11.INJECT1_0 = "NO";
    defparam add_1795_11.INJECT1_1 = "NO";
    LUT4 i22039_4_lut_rep_336 (.A(n31593), .B(count[13]), .C(count[12]), 
         .D(n29377), .Z(n31480)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i22039_4_lut_rep_336.init = 16'heaaa;
    IFS1P3DX latched_in_45 (.D(rc_ch8_c), .SP(n33387), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1246));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1246), .SP(n33387), .CK(debug_c_c), .Q(n1234));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_356_4_lut (.A(count[12]), .B(n31593), .C(count[13]), 
         .D(n31543), .Z(n31500)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_356_4_lut.init = 16'hfffe;
    CCU2D add_1795_9 (.A0(count[7]), .B0(n31602), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n31602), .C1(GND_net), .D1(GND_net), .CIN(n26459), 
          .COUT(n26460), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1795_9.INIT0 = 16'hd222;
    defparam add_1795_9.INIT1 = 16'hd222;
    defparam add_1795_9.INJECT1_0 = "NO";
    defparam add_1795_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(count[4]), .B(n31543), .C(n29253), .D(n4), .Z(n29377)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hfcec;
    CCU2D add_1795_7 (.A0(count[5]), .B0(n31602), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n31602), .C1(GND_net), .D1(GND_net), .CIN(n26458), 
          .COUT(n26459), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1795_7.INIT0 = 16'hd222;
    defparam add_1795_7.INIT1 = 16'hd222;
    defparam add_1795_7.INJECT1_0 = "NO";
    defparam add_1795_7.INJECT1_1 = "NO";
    CCU2D add_1795_5 (.A0(count[3]), .B0(n31602), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n31602), .C1(GND_net), .D1(GND_net), .CIN(n26457), 
          .COUT(n26458), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1795_5.INIT0 = 16'hd222;
    defparam add_1795_5.INIT1 = 16'hd222;
    defparam add_1795_5.INJECT1_0 = "NO";
    defparam add_1795_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_324_3_lut_4_lut (.A(count[9]), .B(n31594), .C(count[8]), 
         .D(n31531), .Z(n31468)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_324_3_lut_4_lut.init = 16'hfffe;
    CCU2D add_1795_3 (.A0(count[1]), .B0(n31602), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n31602), .C1(GND_net), .D1(GND_net), .CIN(n26456), 
          .COUT(n26457), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1795_3.INIT0 = 16'hd222;
    defparam add_1795_3.INIT1 = 16'hd222;
    defparam add_1795_3.INJECT1_0 = "NO";
    defparam add_1795_3.INJECT1_1 = "NO";
    CCU2D add_1795_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29400), .B1(n1246), .C1(count[0]), .D1(n1234), .COUT(n26456), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1795_1.INIT0 = 16'hF000;
    defparam add_1795_1.INIT1 = 16'ha565;
    defparam add_1795_1.INJECT1_0 = "NO";
    defparam add_1795_1.INJECT1_1 = "NO";
    LUT4 i21_3_lut_4_lut (.A(n31531), .B(n31543), .C(n27756), .D(n29314), 
         .Z(n54)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;
    defparam i21_3_lut_4_lut.init = 16'h0f0e;
    LUT4 i22358_4_lut (.A(n54), .B(n29554), .C(n23), .D(n10), .Z(n29818)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i22358_4_lut.init = 16'h3332;
    LUT4 i3_4_lut (.A(n31593), .B(n28997), .C(n31594), .D(n33386), .Z(n17066)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut.init = 16'h0400;
    LUT4 i4_4_lut (.A(count[13]), .B(n24), .C(count[12]), .D(n29554), 
         .Z(n28997)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0004;
    LUT4 i31_3_lut (.A(n29314), .B(n27592), .C(count[9]), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i31_3_lut.init = 16'h3a3a;
    LUT4 i1_2_lut (.A(n23), .B(n1138[7]), .Z(n43[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_325 (.A(count[8]), .B(n31500), .C(n31597), .D(n29472), 
         .Z(n23)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;
    defparam i1_4_lut_adj_325.init = 16'h0222;
    LUT4 i1_4_lut_adj_326 (.A(n31597), .B(n31532), .C(count[0]), .D(n29253), 
         .Z(n29314)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_4_lut_adj_326.init = 16'h8000;
    LUT4 i3_4_lut_adj_327 (.A(count[6]), .B(count[8]), .C(count[7]), .D(n29250), 
         .Z(n27592)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_327.init = 16'hfffe;
    LUT4 i1_4_lut_adj_328 (.A(count[2]), .B(n31583), .C(n6), .D(count[0]), 
         .Z(n29250)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_4_lut_adj_328.init = 16'hccc8;
    LUT4 i2_2_lut (.A(count[3]), .B(count[1]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i22000_2_lut (.A(n1234), .B(n1246), .Z(n29554)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i22000_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_rep_439 (.A(count[4]), .B(count[5]), .Z(n31583)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_439.init = 16'h8888;
    LUT4 i3_4_lut_adj_329 (.A(count[0]), .B(n31595), .C(n31532), .D(n31597), 
         .Z(n27724)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_329.init = 16'h8000;
    LUT4 i2_4_lut (.A(n31595), .B(count[5]), .C(count[4]), .D(n4_adj_218), 
         .Z(n27395)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_2_lut_rep_388_3_lut (.A(count[4]), .B(count[5]), .C(count[3]), 
         .Z(n31532)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_388_3_lut.init = 16'h8080;
    LUT4 i21920_2_lut_3_lut_4_lut (.A(count[4]), .B(count[5]), .C(n31595), 
         .D(count[3]), .Z(n29472)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i21920_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_adj_330 (.A(n23), .B(n1138[6]), .Z(n43[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_330.init = 16'h8888;
    LUT4 i1_2_lut_adj_331 (.A(n23), .B(n1138[5]), .Z(n43[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_331.init = 16'h8888;
    LUT4 i1_2_lut_adj_332 (.A(n23), .B(n1138[4]), .Z(n43[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_332.init = 16'h8888;
    LUT4 i1_2_lut_adj_333 (.A(n23), .B(n1138[3]), .Z(n43[3])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_333.init = 16'h8888;
    LUT4 i1_2_lut_adj_334 (.A(n23), .B(n1138[2]), .Z(n43[2])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_334.init = 16'h8888;
    LUT4 i22462_3_lut_3_lut_4_lut (.A(n27395), .B(n31468), .C(n27756), 
         .D(n31480), .Z(n29401)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i22462_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i1_2_lut_adj_335 (.A(n23), .B(n1138[1]), .Z(n43[1])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_335.init = 16'h8888;
    LUT4 i1_2_lut_rep_449 (.A(count[15]), .B(count[14]), .Z(n31593)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_449.init = 16'heeee;
    LUT4 i2_3_lut_rep_387_4_lut (.A(count[15]), .B(count[14]), .C(count[13]), 
         .D(count[12]), .Z(n31531)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_387_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_450 (.A(count[11]), .B(count[10]), .Z(n31594)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_450.init = 16'heeee;
    LUT4 i1_2_lut_rep_399_3_lut (.A(count[11]), .B(count[10]), .C(count[9]), 
         .Z(n31543)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_399_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_451 (.A(count[6]), .B(count[7]), .Z(n31595)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_451.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), .Z(n29253)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_453 (.A(count[2]), .B(count[1]), .Z(n31597)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_453.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_336 (.A(count[2]), .B(count[1]), .C(count[3]), 
         .Z(n4_adj_218)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_adj_336.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[2]), .B(count[1]), .C(count[5]), .D(count[3]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i5_2_lut_rep_458 (.A(n1234), .B(n1246), .Z(n31602)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_458.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_337 (.A(n1234), .B(n1246), .C(n31480), .Z(n29400)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut_adj_337.init = 16'hf4f4;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n13957), .PD(n17066), .CK(debug_c_c), 
            .Q(\register[6] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n13957), .PD(n17066), .CK(debug_c_c), 
            .Q(\register[6] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n13957), .PD(n17066), .CK(debug_c_c), 
            .Q(\register[6] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n13957), .PD(n17066), .CK(debug_c_c), 
            .Q(\register[6] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n13957), .PD(n17066), .CK(debug_c_c), 
            .Q(\register[6] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n13957), .PD(n17066), .CK(debug_c_c), 
            .Q(\register[6] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n13957), .PD(n17066), .CK(debug_c_c), 
            .Q(\register[6] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D add_1795_17 (.A0(count[15]), .B0(n31602), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26463), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1795_17.INIT0 = 16'hd222;
    defparam add_1795_17.INIT1 = 16'h0000;
    defparam add_1795_17.INJECT1_0 = "NO";
    defparam add_1795_17.INJECT1_1 = "NO";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n13957), .PD(n17066), .CK(debug_c_c), 
            .Q(\register[6] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    FD1P3IX valid_48 (.D(n29401), .SP(n27564), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1240));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_338 (.A(n23), .B(n1138[0]), .Z(n43[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_338.init = 16'h8888;
    CCU2D add_1795_15 (.A0(count[13]), .B0(n31602), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n31602), .C1(GND_net), .D1(GND_net), .CIN(n26462), 
          .COUT(n26463), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1795_15.INIT0 = 16'hd222;
    defparam add_1795_15.INIT1 = 16'hd222;
    defparam add_1795_15.INJECT1_0 = "NO";
    defparam add_1795_15.INJECT1_1 = "NO";
    CCU2D add_1795_13 (.A0(count[11]), .B0(n31602), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n31602), .C1(GND_net), .D1(GND_net), .CIN(n26461), 
          .COUT(n26462), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1795_13.INIT0 = 16'hd222;
    defparam add_1795_13.INIT1 = 16'hd222;
    defparam add_1795_13.INJECT1_0 = "NO";
    defparam add_1795_13.INJECT1_1 = "NO";
    LUT4 i22324_4_lut (.A(n28988), .B(n31602), .C(n31480), .D(n29554), 
         .Z(n29784)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i22324_4_lut.init = 16'h3031;
    LUT4 i3_4_lut_adj_339 (.A(n31468), .B(n31594), .C(n29562), .D(n29638), 
         .Z(n28988)) /* synthesis lut_function=(!(A (B+(D))+!A (B+((D)+!C)))) */ ;
    defparam i3_4_lut_adj_339.init = 16'h0032;
    LUT4 i1_2_lut_adj_340 (.A(n27724), .B(n27395), .Z(n29562)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_340.init = 16'h8888;
    LUT4 i22079_4_lut (.A(n54), .B(n31531), .C(n23), .D(n31467), .Z(n29638)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22079_4_lut.init = 16'hfffe;
    CCU2D sub_79_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26735), 
          .S0(n1138[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_79_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_79_add_2_9.INIT1 = 16'h0000;
    defparam sub_79_add_2_9.INJECT1_0 = "NO";
    defparam sub_79_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_79_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26734), 
          .COUT(n26735), .S0(n1138[5]), .S1(n1138[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_79_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_79_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_79_add_2_7.INJECT1_0 = "NO";
    defparam sub_79_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_79_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26733), 
          .COUT(n26734), .S0(n1138[3]), .S1(n1138[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_79_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_79_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_79_add_2_5.INJECT1_0 = "NO";
    defparam sub_79_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_79_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26732), 
          .COUT(n26733), .S0(n1138[1]), .S1(n1138[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_79_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_79_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_79_add_2_3.INJECT1_0 = "NO";
    defparam sub_79_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_79_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26732), 
          .S1(n1138[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_79_add_2_1.INIT0 = 16'hF000;
    defparam sub_79_add_2_1.INIT1 = 16'h5555;
    defparam sub_79_add_2_1.INJECT1_0 = "NO";
    defparam sub_79_add_2_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U1
//

module PWMReceiver_U1 (\register[5] , debug_c_c, n33386, n33387, rc_ch7_c, 
            GND_net, n33388, n1225, n27543, n29827) /* synthesis syn_module_defined=1 */ ;
    output [7:0]\register[5] ;
    input debug_c_c;
    input n33386;
    input n33387;
    input rc_ch7_c;
    input GND_net;
    input n33388;
    output n1225;
    input n27543;
    output n29827;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n14451, n16852;
    wire [7:0]n43;
    
    wire n31606, n29608, n54;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n79, n31608, n4, n27303, n1231, n1219, n31604, n31509, 
        n31511, n29281, n13768, n31485, n31607, n31510, n31548, 
        n27715, n31605, n29406, n27589, n31484, n31547, n31453, 
        n29580, n31546, n31452, n29407;
    wire [15:0]n116;
    
    wire n26471, n26470, n26469, n26468, n26467, n13402, n26466, 
        n4_adj_217, n26465, n31486, n26464, n27542, n29630, n26739;
    wire [7:0]n1129;
    
    wire n27615, n6, n26738, n26737, n26736, n28967, n24;
    
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14451), .PD(n16852), .CK(debug_c_c), 
            .Q(\register[5] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i22336_4_lut_4_lut (.A(n31606), .B(n29608), .C(n33386), .D(n54), 
         .Z(n14451)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i22336_4_lut_4_lut.init = 16'h5040;
    LUT4 i1_2_lut (.A(count[5]), .B(count[4]), .Z(n79)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i2_4_lut (.A(n31608), .B(count[4]), .C(count[5]), .D(n4), .Z(n27303)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'ha080;
    IFS1P3DX latched_in_45 (.D(rc_ch7_c), .SP(n33387), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1231));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1231), .SP(n33387), .CK(debug_c_c), .Q(n1219));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i21_3_lut_4_lut (.A(n31604), .B(n31509), .C(n31511), .D(n29281), 
         .Z(n54)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i21_3_lut_4_lut.init = 16'h1110;
    LUT4 i1_2_lut_rep_341_3_lut_4_lut (.A(count[9]), .B(n31604), .C(count[8]), 
         .D(n13768), .Z(n31485)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_341_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_366_4_lut (.A(count[3]), .B(n31607), .C(n79), .D(n31608), 
         .Z(n31510)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_366_4_lut.init = 16'h8000;
    LUT4 i5_2_lut_rep_404 (.A(n1219), .B(n1231), .Z(n31548)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_404.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n1219), .B(n1231), .C(n27715), .D(n31605), 
         .Z(n29406)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff4;
    LUT4 i1_3_lut_rep_365 (.A(n27589), .B(n13768), .C(count[9]), .Z(n31509)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_3_lut_rep_365.init = 16'hecec;
    LUT4 i2_2_lut_rep_340_4_lut (.A(n27589), .B(n13768), .C(count[9]), 
         .D(n31604), .Z(n31484)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i2_2_lut_rep_340_4_lut.init = 16'hffec;
    LUT4 i1_3_lut_rep_309_4_lut (.A(n31608), .B(n31547), .C(n31511), .D(count[8]), 
         .Z(n31453)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_3_lut_rep_309_4_lut.init = 16'h0700;
    LUT4 i1_2_lut_3_lut_4_lut_adj_312 (.A(n31608), .B(n31547), .C(n27303), 
         .D(count[0]), .Z(n29580)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_4_lut_adj_312.init = 16'h8000;
    LUT4 i1_2_lut_rep_308_3_lut_4_lut (.A(n13768), .B(n31546), .C(n27303), 
         .D(count[8]), .Z(n31452)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_308_3_lut_4_lut.init = 16'hfffe;
    LUT4 i22460_3_lut_3_lut_4_lut (.A(n31605), .B(n27715), .C(n31452), 
         .D(n31484), .Z(n29407)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i22460_3_lut_3_lut_4_lut.init = 16'h0010;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    CCU2D add_1791_17 (.A0(count[15]), .B0(n31548), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26471), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1791_17.INIT0 = 16'hd222;
    defparam add_1791_17.INIT1 = 16'h0000;
    defparam add_1791_17.INJECT1_0 = "NO";
    defparam add_1791_17.INJECT1_1 = "NO";
    CCU2D add_1791_15 (.A0(count[13]), .B0(n31548), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n31548), .C1(GND_net), .D1(GND_net), .CIN(n26470), 
          .COUT(n26471), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1791_15.INIT0 = 16'hd222;
    defparam add_1791_15.INIT1 = 16'hd222;
    defparam add_1791_15.INJECT1_0 = "NO";
    defparam add_1791_15.INJECT1_1 = "NO";
    CCU2D add_1791_13 (.A0(count[11]), .B0(n31548), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n31548), .C1(GND_net), .D1(GND_net), .CIN(n26469), 
          .COUT(n26470), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1791_13.INIT0 = 16'hd222;
    defparam add_1791_13.INIT1 = 16'hd222;
    defparam add_1791_13.INJECT1_0 = "NO";
    defparam add_1791_13.INJECT1_1 = "NO";
    CCU2D add_1791_11 (.A0(count[9]), .B0(n31548), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n31548), .C1(GND_net), .D1(GND_net), .CIN(n26468), 
          .COUT(n26469), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1791_11.INIT0 = 16'hd222;
    defparam add_1791_11.INIT1 = 16'hd222;
    defparam add_1791_11.INJECT1_0 = "NO";
    defparam add_1791_11.INJECT1_1 = "NO";
    CCU2D add_1791_9 (.A0(count[7]), .B0(n31548), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n31548), .C1(GND_net), .D1(GND_net), .CIN(n26467), 
          .COUT(n26468), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1791_9.INIT0 = 16'hd222;
    defparam add_1791_9.INIT1 = 16'hd222;
    defparam add_1791_9.INJECT1_0 = "NO";
    defparam add_1791_9.INJECT1_1 = "NO";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14451), .PD(n16852), .CK(debug_c_c), 
            .Q(\register[5] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14451), .PD(n16852), .CK(debug_c_c), 
            .Q(\register[5] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14451), .PD(n16852), .CK(debug_c_c), 
            .Q(\register[5] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_313 (.A(count[13]), .B(count[12]), .C(n13402), .D(n31546), 
         .Z(n27715)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_313.init = 16'h8880;
    CCU2D add_1791_7 (.A0(count[5]), .B0(n31548), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n31548), .C1(GND_net), .D1(GND_net), .CIN(n26466), 
          .COUT(n26467), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1791_7.INIT0 = 16'hd222;
    defparam add_1791_7.INIT1 = 16'hd222;
    defparam add_1791_7.INJECT1_0 = "NO";
    defparam add_1791_7.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_314 (.A(n31608), .B(count[5]), .C(count[8]), .D(n4_adj_217), 
         .Z(n13402)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_314.init = 16'ha080;
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14451), .PD(n16852), .CK(debug_c_c), 
            .Q(\register[5] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14451), .PD(n16852), .CK(debug_c_c), 
            .Q(\register[5] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14451), .PD(n16852), .CK(debug_c_c), 
            .Q(\register[5] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14451), .PD(n16852), .CK(debug_c_c), 
            .Q(\register[5] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_460 (.A(count[11]), .B(count[10]), .Z(n31604)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_460.init = 16'heeee;
    LUT4 i1_2_lut_rep_402_3_lut (.A(count[11]), .B(count[10]), .C(count[9]), 
         .Z(n31546)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_402_3_lut.init = 16'hfefe;
    CCU2D add_1791_5 (.A0(count[3]), .B0(n31548), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n31548), .C1(GND_net), .D1(GND_net), .CIN(n26465), 
          .COUT(n26466), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1791_5.INIT0 = 16'hd222;
    defparam add_1791_5.INIT1 = 16'hd222;
    defparam add_1791_5.INJECT1_0 = "NO";
    defparam add_1791_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_367_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(n13768), 
         .D(count[9]), .Z(n31511)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_367_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_461 (.A(count[15]), .B(count[14]), .Z(n31605)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_461.init = 16'heeee;
    LUT4 i2_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(count[13]), 
         .D(count[12]), .Z(n13768)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21912_2_lut_rep_462 (.A(n1219), .B(n1231), .Z(n31606)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i21912_2_lut_rep_462.init = 16'hdddd;
    LUT4 i3069_2_lut_rep_463 (.A(count[1]), .B(count[2]), .Z(n31607)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3069_2_lut_rep_463.init = 16'h8888;
    LUT4 i3_3_lut_rep_403_4_lut (.A(count[1]), .B(count[2]), .C(n79), 
         .D(count[3]), .Z(n31547)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_3_lut_rep_403_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut (.A(count[1]), .B(count[2]), .C(count[3]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[1]), .B(count[2]), .C(count[3]), .D(count[4]), 
         .Z(n4_adj_217)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i1_2_lut_rep_464 (.A(count[7]), .B(count[6]), .Z(n31608)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_464.init = 16'h8888;
    LUT4 i1_2_lut_rep_342_3_lut_4_lut (.A(count[7]), .B(count[6]), .C(count[0]), 
         .D(n31547), .Z(n31486)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_342_3_lut_4_lut.init = 16'h8000;
    CCU2D add_1791_3 (.A0(count[1]), .B0(n31548), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n31548), .C1(GND_net), .D1(GND_net), .CIN(n26464), 
          .COUT(n26465), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1791_3.INIT0 = 16'hd222;
    defparam add_1791_3.INIT1 = 16'hd222;
    defparam add_1791_3.INJECT1_0 = "NO";
    defparam add_1791_3.INJECT1_1 = "NO";
    CCU2D add_1791_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29406), .B1(n1231), .C1(count[0]), .D1(n1219), .COUT(n26464), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1791_1.INIT0 = 16'hF000;
    defparam add_1791_1.INIT1 = 16'ha565;
    defparam add_1791_1.INJECT1_0 = "NO";
    defparam add_1791_1.INJECT1_1 = "NO";
    FD1P3IX valid_48 (.D(n29407), .SP(n27543), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1225));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i22367_4_lut (.A(n31605), .B(n31548), .C(n27715), .D(n27542), 
         .Z(n29827)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i22367_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n31485), .B(n31606), .C(n29630), .D(n29580), .Z(n27542)) /* synthesis lut_function=(A (B+!(C))+!A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut.init = 16'hcfce;
    LUT4 i22071_4_lut (.A(n31604), .B(n54), .C(n31509), .D(n31453), 
         .Z(n29630)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22071_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_315 (.A(n31547), .B(n31608), .C(count[8]), .D(count[0]), 
         .Z(n29281)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_4_lut_adj_315.init = 16'h8000;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    CCU2D sub_78_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26739), 
          .S0(n1129[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_78_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_78_add_2_9.INIT1 = 16'h0000;
    defparam sub_78_add_2_9.INJECT1_0 = "NO";
    defparam sub_78_add_2_9.INJECT1_1 = "NO";
    LUT4 i3_4_lut (.A(n27615), .B(n6), .C(count[8]), .D(n79), .Z(n27589)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i3_4_lut.init = 16'hfefc;
    CCU2D sub_78_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26738), 
          .COUT(n26739), .S0(n1129[5]), .S1(n1129[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_78_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_78_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_78_add_2_7.INJECT1_0 = "NO";
    defparam sub_78_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_78_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26737), 
          .COUT(n26738), .S0(n1129[3]), .S1(n1129[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_78_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_78_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_78_add_2_5.INJECT1_0 = "NO";
    defparam sub_78_add_2_5.INJECT1_1 = "NO";
    LUT4 i22049_4_lut_4_lut (.A(n27303), .B(n31485), .C(n31486), .D(n31453), 
         .Z(n29608)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (D)) */ ;
    defparam i22049_4_lut_4_lut.init = 16'hff02;
    LUT4 i1_2_lut_4_lut (.A(count[8]), .B(n31510), .C(n31511), .D(n1129[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0200;
    CCU2D sub_78_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26736), 
          .COUT(n26737), .S0(n1129[1]), .S1(n1129[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_78_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_78_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_78_add_2_3.INJECT1_0 = "NO";
    defparam sub_78_add_2_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_316 (.A(count[8]), .B(n31510), .C(n31511), 
         .D(n1129[1]), .Z(n43[1])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_316.init = 16'h0200;
    LUT4 i1_2_lut_4_lut_adj_317 (.A(count[8]), .B(n31510), .C(n31511), 
         .D(n1129[4]), .Z(n43[4])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_317.init = 16'h0200;
    LUT4 i1_2_lut_4_lut_adj_318 (.A(count[8]), .B(n31510), .C(n31511), 
         .D(n1129[5]), .Z(n43[5])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_318.init = 16'h0200;
    CCU2D sub_78_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26736), 
          .S1(n1129[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_78_add_2_1.INIT0 = 16'hF000;
    defparam sub_78_add_2_1.INIT1 = 16'h5555;
    defparam sub_78_add_2_1.INJECT1_0 = "NO";
    defparam sub_78_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_319 (.A(count[8]), .B(n31510), .C(n31511), 
         .D(n1129[6]), .Z(n43[6])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_319.init = 16'h0200;
    LUT4 i1_2_lut_4_lut_adj_320 (.A(count[8]), .B(n31510), .C(n31511), 
         .D(n1129[7]), .Z(n43[7])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_320.init = 16'h0200;
    LUT4 i1_2_lut_4_lut_adj_321 (.A(count[8]), .B(n31510), .C(n31511), 
         .D(n1129[0]), .Z(n43[0])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_321.init = 16'h0200;
    LUT4 i3_4_lut_adj_322 (.A(count[0]), .B(count[1]), .C(count[3]), .D(count[2]), 
         .Z(n27615)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_322.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_323 (.A(count[8]), .B(n31510), .C(n31511), 
         .D(n1129[2]), .Z(n43[2])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_323.init = 16'h0200;
    LUT4 i2_2_lut (.A(count[6]), .B(count[7]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_324 (.A(n31605), .B(n28967), .C(n31604), .D(n33386), 
         .Z(n16852)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_324.init = 16'h0400;
    LUT4 i4_4_lut (.A(count[13]), .B(n24), .C(count[12]), .D(n31606), 
         .Z(n28967)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0004;
    LUT4 i31_3_lut (.A(n29281), .B(n27589), .C(count[9]), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i31_3_lut.init = 16'h3a3a;
    
endmodule
//
// Verilog Description of module PWMReceiver_U2
//

module PWMReceiver_U2 (n33386, debug_c_c, n33387, rc_ch4_c, GND_net, 
            n33388, \register[4] , n1210, n27550, n29838) /* synthesis syn_module_defined=1 */ ;
    input n33386;
    input debug_c_c;
    input n33387;
    input rc_ch4_c;
    input GND_net;
    input n33388;
    output [7:0]\register[4] ;
    output n1210;
    input n27550;
    output n29838;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n31559, n31517, n29291, n31558, n124, n31489, n31555, 
        n4, n31433, n14491, n31557, n27645, n31434, n22311, n29316, 
        n1216, n1204, n31490, n31456, n5, n27366, n31455, n29305, 
        n13677, n5_adj_212, n29317, n4_adj_213, n4_adj_214, n31516, 
        n31560, n29644, n31564, n103, n26479;
    wire [15:0]n116;
    
    wire n26478, n26477, n26476, n152, n154, n16891;
    wire [7:0]n43;
    
    wire n26475, n26474, n26473, n26472, n6, n29577, n4_adj_216;
    wire [7:0]n1120;
    
    wire n11, n8, n27548, n26743, n26742, n26741, n26740;
    
    LUT4 i1_3_lut_4_lut (.A(count[8]), .B(n31559), .C(count[0]), .D(n31517), 
         .Z(n29291)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_345_4_lut (.A(count[3]), .B(n31558), .C(n124), .D(n31559), 
         .Z(n31489)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_345_4_lut.init = 16'h8000;
    LUT4 i22488_4_lut_4_lut (.A(n31555), .B(n4), .C(n33386), .D(n31433), 
         .Z(n14491)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i22488_4_lut_4_lut.init = 16'h5010;
    LUT4 i22455_3_lut_3_lut_4_lut (.A(n31557), .B(n27645), .C(n31434), 
         .D(n22311), .Z(n29316)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i22455_3_lut_3_lut_4_lut.init = 16'h0010;
    IFS1P3DX latched_in_45 (.D(rc_ch4_c), .SP(n33387), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1216));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1216), .SP(n33387), .CK(debug_c_c), .Q(n1204));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut (.A(n29291), .B(n22311), .C(n31490), .D(n31456), 
         .Z(n5)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i1_2_lut_4_lut.init = 16'hcd00;
    LUT4 i1_4_lut_4_lut (.A(n27366), .B(n31455), .C(n29305), .D(n31456), 
         .Z(n4)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i1_4_lut_4_lut.init = 16'hfd00;
    LUT4 i1_3_lut_rep_312_4_lut (.A(n31559), .B(n31517), .C(count[8]), 
         .D(n31490), .Z(n31456)) /* synthesis lut_function=(A (B+((D)+!C))+!A ((D)+!C)) */ ;
    defparam i1_3_lut_rep_312_4_lut.init = 16'hff8f;
    LUT4 i1_2_lut_rep_346 (.A(count[9]), .B(n13677), .Z(n31490)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_346.init = 16'heeee;
    LUT4 i1_2_lut_rep_311_3_lut (.A(count[9]), .B(n13677), .C(count[8]), 
         .Z(n31455)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_311_3_lut.init = 16'hfefe;
    LUT4 i21_3_lut_rep_289_4_lut (.A(count[9]), .B(n13677), .C(n22311), 
         .D(n29291), .Z(n31433)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i21_3_lut_rep_289_4_lut.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_290_3_lut_4_lut (.A(count[9]), .B(n13677), .C(n27366), 
         .D(count[8]), .Z(n31434)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_290_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_411 (.A(n1216), .B(n1204), .Z(n31555)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_411.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_413 (.A(count[15]), .B(count[14]), .Z(n31557)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_413.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(n5_adj_212), 
         .D(n27645), .Z(n29317)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_414 (.A(count[2]), .B(count[1]), .Z(n31558)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_414.init = 16'h8888;
    LUT4 i1_3_lut_rep_373_4_lut (.A(count[2]), .B(count[1]), .C(n124), 
         .D(count[3]), .Z(n31517)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_3_lut_rep_373_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[4]), .Z(n4_adj_213)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut_adj_305 (.A(count[2]), .B(count[1]), .C(count[5]), 
         .D(count[3]), .Z(n4_adj_214)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut_adj_305.init = 16'hf8f0;
    LUT4 i1_2_lut_rep_415 (.A(count[7]), .B(count[6]), .Z(n31559)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_415.init = 16'h8888;
    LUT4 i1_2_lut_rep_372_3_lut (.A(count[7]), .B(count[6]), .C(count[8]), 
         .Z(n31516)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_372_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_306 (.A(count[7]), .B(count[6]), .C(count[0]), 
         .D(n31517), .Z(n29305)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_4_lut_adj_306.init = 16'h8000;
    LUT4 i21936_2_lut_rep_416 (.A(count[11]), .B(count[10]), .Z(n31560)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21936_2_lut_rep_416.init = 16'heeee;
    LUT4 i22085_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(count[13]), 
         .D(count[12]), .Z(n29644)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22085_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_420 (.A(count[7]), .B(count[6]), .C(count[8]), .Z(n31564)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_420.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_307 (.A(count[7]), .B(count[6]), .C(count[8]), 
         .D(n124), .Z(n103)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_307.init = 16'hfffe;
    CCU2D add_1787_17 (.A0(count[15]), .B0(n5_adj_212), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26479), .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1787_17.INIT0 = 16'hd222;
    defparam add_1787_17.INIT1 = 16'h0000;
    defparam add_1787_17.INJECT1_0 = "NO";
    defparam add_1787_17.INJECT1_1 = "NO";
    CCU2D add_1787_15 (.A0(count[13]), .B0(n5_adj_212), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n5_adj_212), .C1(GND_net), 
          .D1(GND_net), .CIN(n26478), .COUT(n26479), .S0(n116[13]), 
          .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1787_15.INIT0 = 16'hd222;
    defparam add_1787_15.INIT1 = 16'hd222;
    defparam add_1787_15.INJECT1_0 = "NO";
    defparam add_1787_15.INJECT1_1 = "NO";
    CCU2D add_1787_13 (.A0(count[11]), .B0(n5_adj_212), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n5_adj_212), .C1(GND_net), 
          .D1(GND_net), .CIN(n26477), .COUT(n26478), .S0(n116[11]), 
          .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1787_13.INIT0 = 16'hd222;
    defparam add_1787_13.INIT1 = 16'hd222;
    defparam add_1787_13.INJECT1_0 = "NO";
    defparam add_1787_13.INJECT1_1 = "NO";
    CCU2D add_1787_11 (.A0(count[9]), .B0(n5_adj_212), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5_adj_212), .C1(GND_net), .D1(GND_net), 
          .CIN(n26476), .COUT(n26477), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1787_11.INIT0 = 16'hd222;
    defparam add_1787_11.INIT1 = 16'hd222;
    defparam add_1787_11.INJECT1_0 = "NO";
    defparam add_1787_11.INJECT1_1 = "NO";
    PFUMX i14066 (.BLUT(n152), .ALUT(n103), .C0(count[3]), .Z(n154));
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14491), .PD(n16891), .CK(debug_c_c), 
            .Q(\register[4] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14491), .PD(n16891), .CK(debug_c_c), 
            .Q(\register[4] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    CCU2D add_1787_9 (.A0(count[7]), .B0(n5_adj_212), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5_adj_212), .C1(GND_net), .D1(GND_net), 
          .CIN(n26475), .COUT(n26476), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1787_9.INIT0 = 16'hd222;
    defparam add_1787_9.INIT1 = 16'hd222;
    defparam add_1787_9.INJECT1_0 = "NO";
    defparam add_1787_9.INJECT1_1 = "NO";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14491), .PD(n16891), .CK(debug_c_c), 
            .Q(\register[4] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14491), .PD(n16891), .CK(debug_c_c), 
            .Q(\register[4] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14491), .PD(n16891), .CK(debug_c_c), 
            .Q(\register[4] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14491), .PD(n16891), .CK(debug_c_c), 
            .Q(\register[4] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14491), .PD(n16891), .CK(debug_c_c), 
            .Q(\register[4] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D add_1787_7 (.A0(count[5]), .B0(n5_adj_212), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5_adj_212), .C1(GND_net), .D1(GND_net), 
          .CIN(n26474), .COUT(n26475), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1787_7.INIT0 = 16'hd222;
    defparam add_1787_7.INIT1 = 16'hd222;
    defparam add_1787_7.INJECT1_0 = "NO";
    defparam add_1787_7.INJECT1_1 = "NO";
    CCU2D add_1787_5 (.A0(count[3]), .B0(n5_adj_212), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5_adj_212), .C1(GND_net), .D1(GND_net), 
          .CIN(n26473), .COUT(n26474), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1787_5.INIT0 = 16'hd222;
    defparam add_1787_5.INIT1 = 16'hd222;
    defparam add_1787_5.INJECT1_0 = "NO";
    defparam add_1787_5.INJECT1_1 = "NO";
    CCU2D add_1787_3 (.A0(count[1]), .B0(n5_adj_212), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5_adj_212), .C1(GND_net), .D1(GND_net), 
          .CIN(n26472), .COUT(n26473), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1787_3.INIT0 = 16'hd222;
    defparam add_1787_3.INIT1 = 16'hd222;
    defparam add_1787_3.INJECT1_0 = "NO";
    defparam add_1787_3.INJECT1_1 = "NO";
    CCU2D add_1787_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29317), .B1(n1216), .C1(count[0]), .D1(n1204), .COUT(n26472), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1787_1.INIT0 = 16'hF000;
    defparam add_1787_1.INIT1 = 16'ha565;
    defparam add_1787_1.INJECT1_0 = "NO";
    defparam add_1787_1.INJECT1_1 = "NO";
    LUT4 i23_4_lut (.A(n31564), .B(count[2]), .C(n124), .D(n6), .Z(n152)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'hfaea;
    LUT4 i2_2_lut (.A(count[1]), .B(count[0]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1_2_lut (.A(count[4]), .B(count[5]), .Z(n124)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i22020_3_lut_4_lut (.A(count[8]), .B(n31490), .C(n27366), .D(n29305), 
         .Z(n29577)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i22020_3_lut_4_lut.init = 16'hfeee;
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n31560), .D(n4_adj_216), 
         .Z(n27645)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_4_lut (.A(count[9]), .B(count[4]), .C(n31516), .D(n4_adj_214), 
         .Z(n4_adj_216)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'hfaea;
    LUT4 i15417_2_lut_4_lut (.A(n31490), .B(count[8]), .C(n31489), .D(n1120[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15417_2_lut_4_lut.init = 16'h0400;
    LUT4 i2_4_lut_adj_308 (.A(n33386), .B(n31557), .C(n11), .D(n29644), 
         .Z(n16891)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut_adj_308.init = 16'h0020;
    LUT4 i15416_2_lut_4_lut (.A(n31490), .B(count[8]), .C(n31489), .D(n1120[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15416_2_lut_4_lut.init = 16'h0400;
    LUT4 i15415_2_lut_4_lut (.A(n31490), .B(count[8]), .C(n31489), .D(n1120[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15415_2_lut_4_lut.init = 16'h0400;
    LUT4 i4_4_lut (.A(n29291), .B(n8), .C(n154), .D(count[9]), .Z(n11)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A ((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i4_4_lut.init = 16'h0c88;
    FD1P3IX valid_48 (.D(n29316), .SP(n27550), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1210));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i22378_4_lut (.A(n31557), .B(n5_adj_212), .C(n27645), .D(n27548), 
         .Z(n29838)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i22378_4_lut.init = 16'h3233;
    LUT4 i1_4_lut_adj_309 (.A(n5), .B(n31555), .C(n29577), .D(n22311), 
         .Z(n27548)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut_adj_309.init = 16'hccec;
    LUT4 i15414_2_lut_4_lut (.A(n31490), .B(count[8]), .C(n31489), .D(n1120[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15414_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_adj_310 (.A(n1204), .B(n1216), .Z(n8)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_adj_310.init = 16'h2222;
    LUT4 i15413_2_lut_4_lut (.A(n31490), .B(count[8]), .C(n31489), .D(n1120[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15413_2_lut_4_lut.init = 16'h0400;
    LUT4 i15412_2_lut_4_lut (.A(n31490), .B(count[8]), .C(n31489), .D(n1120[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15412_2_lut_4_lut.init = 16'h0400;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14491), .PD(n16891), .CK(debug_c_c), 
            .Q(\register[4] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i15411_2_lut_4_lut (.A(n31490), .B(count[8]), .C(n31489), .D(n1120[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15411_2_lut_4_lut.init = 16'h0400;
    LUT4 i15197_2_lut_4_lut (.A(n31490), .B(count[8]), .C(n31489), .D(n1120[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15197_2_lut_4_lut.init = 16'h0400;
    CCU2D sub_77_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26743), 
          .S0(n1120[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_77_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_77_add_2_9.INIT1 = 16'h0000;
    defparam sub_77_add_2_9.INJECT1_0 = "NO";
    defparam sub_77_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_77_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26742), 
          .COUT(n26743), .S0(n1120[5]), .S1(n1120[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_77_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_77_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_77_add_2_7.INJECT1_0 = "NO";
    defparam sub_77_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_77_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26741), 
          .COUT(n26742), .S0(n1120[3]), .S1(n1120[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_77_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_77_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_77_add_2_5.INJECT1_0 = "NO";
    defparam sub_77_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_77_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26740), 
          .COUT(n26741), .S0(n1120[1]), .S1(n1120[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_77_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_77_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_77_add_2_3.INJECT1_0 = "NO";
    defparam sub_77_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_77_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26740), 
          .S1(n1120[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_77_add_2_1.INIT0 = 16'hF000;
    defparam sub_77_add_2_1.INIT1 = 16'h5555;
    defparam sub_77_add_2_1.INJECT1_0 = "NO";
    defparam sub_77_add_2_1.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_311 (.A(n31559), .B(count[5]), .C(count[3]), .D(n4_adj_213), 
         .Z(n27366)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_311.init = 16'h8880;
    LUT4 i3_4_lut (.A(count[12]), .B(count[13]), .C(n31557), .D(n31560), 
         .Z(n13677)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(n1204), .B(n1216), .Z(n5_adj_212)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i15575_3_lut (.A(count[9]), .B(n13677), .C(n154), .Z(n22311)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i15575_3_lut.init = 16'hecec;
    
endmodule
//
// Verilog Description of module PWMReceiver_U3
//

module PWMReceiver_U3 (debug_c_c, n33387, rc_ch3_c, GND_net, n33388, 
            \register[3] , n14500, n1195, n27541, n29840, n29530, 
            n29944, n14) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n33387;
    input rc_ch3_c;
    input GND_net;
    input n33388;
    output [7:0]\register[3] ;
    input n14500;
    output n1195;
    input n27541;
    output n29840;
    output n29530;
    output n29944;
    input n14;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n1189, n1201, n5;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n31565, n31572, n31574, n31493, n26487;
    wire [15:0]n116;
    
    wire n26486, n13663, n31492, n31458, n31459, n31522, n29302, 
        n27278, n29592, n31439, n29410, n26485, n154, n26484, 
        n31562, n103, n26483, n5_adj_208, n54, n7, n6, n31525, 
        n4, n4_adj_209, n31575, n27717, n29409, n26482, n26481, 
        n26480;
    wire [7:0]n1111;
    wire [7:0]n43;
    
    wire n16901, n152, n6_adj_210, n27540, n29595, n26747, n26746, 
        n26745, n26744, n29344, n4_adj_211, n10, n29650, n26;
    
    LUT4 i5_2_lut (.A(n1189), .B(n1201), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i3_3_lut_rep_349_4_lut (.A(count[3]), .B(n31565), .C(n31572), 
         .D(n31574), .Z(n31493)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i3_3_lut_rep_349_4_lut.init = 16'h8000;
    IFS1P3DX latched_in_45 (.D(rc_ch3_c), .SP(n33387), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1201));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1201), .SP(n33387), .CK(debug_c_c), .Q(n1189));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    CCU2D add_1783_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26487), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_17.INIT0 = 16'hd222;
    defparam add_1783_17.INIT1 = 16'h0000;
    defparam add_1783_17.INJECT1_0 = "NO";
    defparam add_1783_17.INJECT1_1 = "NO";
    CCU2D add_1783_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26486), 
          .COUT(n26487), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_15.INIT0 = 16'hd222;
    defparam add_1783_15.INIT1 = 16'hd222;
    defparam add_1783_15.INJECT1_0 = "NO";
    defparam add_1783_15.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_348 (.A(count[9]), .B(n13663), .Z(n31492)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_348.init = 16'heeee;
    LUT4 i1_2_lut_rep_314_3_lut (.A(count[9]), .B(n13663), .C(count[8]), 
         .Z(n31458)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_314_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_rep_315_4_lut (.A(count[9]), .B(n13663), .C(n31493), 
         .D(count[8]), .Z(n31459)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i2_3_lut_rep_315_4_lut.init = 16'hfeff;
    LUT4 i1_2_lut_4_lut (.A(n31574), .B(n31572), .C(n31522), .D(count[0]), 
         .Z(n29302)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h8000;
    LUT4 i22453_3_lut_3_lut_4_lut (.A(n27278), .B(n31458), .C(n29592), 
         .D(n31439), .Z(n29410)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i22453_3_lut_3_lut_4_lut.init = 16'h000e;
    CCU2D add_1783_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26485), 
          .COUT(n26486), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_13.INIT0 = 16'hd222;
    defparam add_1783_13.INIT1 = 16'hd222;
    defparam add_1783_13.INJECT1_0 = "NO";
    defparam add_1783_13.INJECT1_1 = "NO";
    LUT4 i22034_3_lut (.A(n13663), .B(count[9]), .C(n154), .Z(n29592)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i22034_3_lut.init = 16'heaea;
    CCU2D add_1783_11 (.A0(count[9]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26484), 
          .COUT(n26485), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_11.INIT0 = 16'hd222;
    defparam add_1783_11.INIT1 = 16'hd222;
    defparam add_1783_11.INJECT1_0 = "NO";
    defparam add_1783_11.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_418 (.A(count[7]), .B(count[6]), .C(count[8]), .Z(n31562)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_418.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_300 (.A(count[7]), .B(count[6]), .C(count[8]), 
         .D(n31565), .Z(n103)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_300.init = 16'hfffe;
    CCU2D add_1783_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26483), 
          .COUT(n26484), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_9.INIT0 = 16'hd222;
    defparam add_1783_9.INIT1 = 16'hd222;
    defparam add_1783_9.INJECT1_0 = "NO";
    defparam add_1783_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_421 (.A(count[4]), .B(count[5]), .Z(n31565)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_421.init = 16'h8888;
    LUT4 i1_2_lut_rep_378_3_lut (.A(count[4]), .B(count[5]), .C(count[3]), 
         .Z(n31522)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_378_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[4]), .B(count[5]), .C(count[0]), 
         .D(count[3]), .Z(n5_adj_208)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_428 (.A(count[7]), .B(count[6]), .Z(n31572)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_428.init = 16'h8888;
    LUT4 i1_2_lut_4_lut_adj_301 (.A(n31492), .B(count[8]), .C(n31493), 
         .D(n54), .Z(n7)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_301.init = 16'h00fb;
    LUT4 i2_2_lut_3_lut_4_lut (.A(count[7]), .B(count[6]), .C(n31574), 
         .D(count[8]), .Z(n6)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_381_3_lut (.A(count[7]), .B(count[6]), .C(count[8]), 
         .Z(n31525)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_381_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_430 (.A(count[2]), .B(count[1]), .Z(n31574)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_430.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[4]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[2]), .B(count[1]), .C(count[5]), .D(count[3]), 
         .Z(n4_adj_209)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_rep_431 (.A(count[15]), .B(count[14]), .Z(n31575)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_431.init = 16'heeee;
    LUT4 i1_2_lut_rep_295_3_lut (.A(count[15]), .B(count[14]), .C(n27717), 
         .Z(n31439)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_295_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_302 (.A(count[15]), .B(count[14]), .C(n5), 
         .D(n27717), .Z(n29409)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_302.init = 16'hfffe;
    CCU2D add_1783_7 (.A0(count[5]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26482), 
          .COUT(n26483), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_7.INIT0 = 16'hd222;
    defparam add_1783_7.INIT1 = 16'hd222;
    defparam add_1783_7.INJECT1_0 = "NO";
    defparam add_1783_7.INJECT1_1 = "NO";
    CCU2D add_1783_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26481), 
          .COUT(n26482), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_5.INIT0 = 16'hd222;
    defparam add_1783_5.INIT1 = 16'hd222;
    defparam add_1783_5.INJECT1_0 = "NO";
    defparam add_1783_5.INJECT1_1 = "NO";
    CCU2D add_1783_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26480), 
          .COUT(n26481), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_3.INIT0 = 16'hd222;
    defparam add_1783_3.INIT1 = 16'hd222;
    defparam add_1783_3.INJECT1_0 = "NO";
    defparam add_1783_3.INJECT1_1 = "NO";
    CCU2D add_1783_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29409), .B1(n1201), .C1(count[0]), .D1(n1189), .COUT(n26480), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_1.INIT0 = 16'hF000;
    defparam add_1783_1.INIT1 = 16'ha565;
    defparam add_1783_1.INJECT1_0 = "NO";
    defparam add_1783_1.INJECT1_1 = "NO";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    LUT4 i15185_2_lut_4_lut (.A(n31492), .B(count[8]), .C(n31493), .D(n1111[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15185_2_lut_4_lut.init = 16'h0400;
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14500), .PD(n16901), .CK(debug_c_c), 
            .Q(\register[3] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    PFUMX i14315 (.BLUT(n152), .ALUT(n103), .C0(count[3]), .Z(n154));
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14500), .PD(n16901), .CK(debug_c_c), 
            .Q(\register[3] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14500), .PD(n16901), .CK(debug_c_c), 
            .Q(\register[3] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14500), .PD(n16901), .CK(debug_c_c), 
            .Q(\register[3] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14500), .PD(n16901), .CK(debug_c_c), 
            .Q(\register[3] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14500), .PD(n16901), .CK(debug_c_c), 
            .Q(\register[3] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14500), .PD(n16901), .CK(debug_c_c), 
            .Q(\register[3] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i23_4_lut (.A(n31562), .B(count[2]), .C(n31565), .D(n6_adj_210), 
         .Z(n152)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'hfaea;
    LUT4 i2_2_lut (.A(count[1]), .B(count[0]), .Z(n6_adj_210)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    FD1P3IX valid_48 (.D(n29410), .SP(n27541), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1195));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i22380_4_lut (.A(n31575), .B(n5), .C(n27717), .D(n27540), .Z(n29840)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i22380_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n29592), .B(n29530), .C(n7), .D(n29595), .Z(n27540)) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hdccc;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14500), .PD(n16901), .CK(debug_c_c), 
            .Q(\register[3] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D sub_76_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26747), 
          .S0(n1111[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_76_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_76_add_2_9.INIT1 = 16'h0000;
    defparam sub_76_add_2_9.INJECT1_0 = "NO";
    defparam sub_76_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_76_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26746), 
          .COUT(n26747), .S0(n1111[5]), .S1(n1111[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_76_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_76_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_76_add_2_7.INJECT1_0 = "NO";
    defparam sub_76_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_76_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26745), 
          .COUT(n26746), .S0(n1111[3]), .S1(n1111[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_76_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_76_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_76_add_2_5.INJECT1_0 = "NO";
    defparam sub_76_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_76_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26744), 
          .COUT(n26745), .S0(n1111[1]), .S1(n1111[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_76_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_76_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_76_add_2_3.INJECT1_0 = "NO";
    defparam sub_76_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_76_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26744), 
          .S1(n1111[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_76_add_2_1.INIT0 = 16'hF000;
    defparam sub_76_add_2_1.INIT1 = 16'h5555;
    defparam sub_76_add_2_1.INJECT1_0 = "NO";
    defparam sub_76_add_2_1.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n29344), .D(n4_adj_211), 
         .Z(n27717)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_4_lut_adj_303 (.A(count[9]), .B(count[4]), .C(n31525), .D(n4_adj_209), 
         .Z(n4_adj_211)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_303.init = 16'hfaea;
    LUT4 i1_2_lut (.A(count[10]), .B(count[11]), .Z(n29344)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n31492), .C(n29302), 
         .D(n27278), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i22036_3_lut_4_lut (.A(count[8]), .B(n31492), .C(n27278), .D(n29302), 
         .Z(n29595)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i22036_3_lut_4_lut.init = 16'hfeee;
    LUT4 i15410_2_lut_4_lut (.A(n31492), .B(count[8]), .C(n31493), .D(n1111[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15410_2_lut_4_lut.init = 16'h0400;
    LUT4 i15409_2_lut_4_lut (.A(n31492), .B(count[8]), .C(n31493), .D(n1111[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15409_2_lut_4_lut.init = 16'h0400;
    LUT4 i15408_2_lut_4_lut (.A(n31492), .B(count[8]), .C(n31493), .D(n1111[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15408_2_lut_4_lut.init = 16'h0400;
    LUT4 i15407_2_lut_4_lut (.A(n31492), .B(count[8]), .C(n31493), .D(n1111[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15407_2_lut_4_lut.init = 16'h0400;
    LUT4 i22484_4_lut (.A(n54), .B(n29530), .C(n31459), .D(n10), .Z(n29944)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i22484_4_lut.init = 16'h3323;
    LUT4 i15406_2_lut_4_lut (.A(n31492), .B(count[8]), .C(n31493), .D(n1111[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15406_2_lut_4_lut.init = 16'h0400;
    LUT4 i8_4_lut (.A(n29650), .B(count[10]), .C(n14), .D(n26), .Z(n16901)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i8_4_lut.init = 16'h1000;
    LUT4 i22091_4_lut (.A(count[12]), .B(count[13]), .C(count[11]), .D(n31575), 
         .Z(n29650)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22091_4_lut.init = 16'hfffe;
    LUT4 i33_4_lut (.A(count[8]), .B(n154), .C(count[9]), .D(n29302), 
         .Z(n26)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i33_4_lut.init = 16'h3a30;
    LUT4 i15405_2_lut_4_lut (.A(n31492), .B(count[8]), .C(n31493), .D(n1111[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15405_2_lut_4_lut.init = 16'h0400;
    LUT4 i15404_2_lut_4_lut (.A(n31492), .B(count[8]), .C(n31493), .D(n1111[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i15404_2_lut_4_lut.init = 16'h0400;
    LUT4 i21976_2_lut (.A(n1189), .B(n1201), .Z(n29530)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i21976_2_lut.init = 16'hdddd;
    LUT4 i2_4_lut_adj_304 (.A(n31572), .B(count[5]), .C(count[3]), .D(n4), 
         .Z(n27278)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_304.init = 16'h8880;
    LUT4 i3_4_lut (.A(count[12]), .B(n31575), .C(count[13]), .D(n29344), 
         .Z(n13663)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(n5_adj_208), .B(n29592), .C(n31492), .D(n6), 
         .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h3230;
    
endmodule
//
// Verilog Description of module PWMReceiver_U4
//

module PWMReceiver_U4 (GND_net, n29832, debug_c_c, n33387, rc_ch2_c, 
            n31412, n33388, \register[2] , n14513, n29847, n1180, 
            n27536, n33386, n31512) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n29832;
    input debug_c_c;
    input n33387;
    input rc_ch2_c;
    input n31412;
    input n33388;
    output [7:0]\register[2] ;
    input n14513;
    output n29847;
    output n1180;
    input n27536;
    input n33386;
    input n31512;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26491;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n31573;
    wire [15:0]n116;
    
    wire n26492, n29351, n27565, n4, n29352, n29187, n26490, n13702, 
        n26489, n26488, n31482, n29397, n1186, n1174, n13631, 
        n31494, n31460, n31495, n22410, n27662, n31437, n129_adj_206, 
        n31461, n29518, n23, n29654, n29398, n31566, n27609, n31570, 
        n31599, n16910;
    wire [7:0]n43;
    
    wire n31438, n18, n29248, n26495, n26751;
    wire [7:0]n1102;
    
    wire n26750, n26749, n26748, n28999, n4_adj_207, n5, n6, n27518, 
        n26494, n26493;
    
    CCU2D add_1779_9 (.A0(count[7]), .B0(n31573), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n31573), .C1(GND_net), .D1(GND_net), .CIN(n26491), 
          .COUT(n26492), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_9.INIT0 = 16'hd222;
    defparam add_1779_9.INIT1 = 16'hd222;
    defparam add_1779_9.INJECT1_0 = "NO";
    defparam add_1779_9.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(n29351), .B(count[9]), .C(n27565), .D(n4), .Z(n29352)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut.init = 16'hfeee;
    LUT4 i2_4_lut_adj_288 (.A(count[1]), .B(count[5]), .C(n29187), .D(count[4]), 
         .Z(n27565)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_288.init = 16'hffec;
    LUT4 i1_2_lut (.A(count[10]), .B(count[11]), .Z(n29351)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_289 (.A(count[3]), .B(count[2]), .Z(n29187)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_adj_289.init = 16'h8888;
    CCU2D add_1779_7 (.A0(count[5]), .B0(n31573), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n31573), .C1(GND_net), .D1(GND_net), .CIN(n26490), 
          .COUT(n26491), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_7.INIT0 = 16'hd222;
    defparam add_1779_7.INIT1 = 16'hd222;
    defparam add_1779_7.INJECT1_0 = "NO";
    defparam add_1779_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_290 (.A(count[15]), .B(count[14]), .Z(n13702)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_290.init = 16'heeee;
    CCU2D add_1779_5 (.A0(count[3]), .B0(n31573), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n31573), .C1(GND_net), .D1(GND_net), .CIN(n26489), 
          .COUT(n26490), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_5.INIT0 = 16'hd222;
    defparam add_1779_5.INIT1 = 16'hd222;
    defparam add_1779_5.INJECT1_0 = "NO";
    defparam add_1779_5.INJECT1_1 = "NO";
    CCU2D add_1779_3 (.A0(count[1]), .B0(n31573), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n31573), .C1(GND_net), .D1(GND_net), .CIN(n26488), 
          .COUT(n26489), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_3.INIT0 = 16'hd222;
    defparam add_1779_3.INIT1 = 16'hd222;
    defparam add_1779_3.INJECT1_0 = "NO";
    defparam add_1779_3.INJECT1_1 = "NO";
    LUT4 i1_4_lut_rep_338 (.A(n13702), .B(count[13]), .C(count[12]), .D(n29352), 
         .Z(n31482)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_rep_338.init = 16'heaaa;
    CCU2D add_1779_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29397), .B1(n1186), .C1(count[0]), .D1(n1174), .COUT(n26488), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_1.INIT0 = 16'hF000;
    defparam add_1779_1.INIT1 = 16'ha565;
    defparam add_1779_1.INJECT1_0 = "NO";
    defparam add_1779_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_350 (.A(count[9]), .B(n13631), .Z(n31494)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_350.init = 16'heeee;
    LUT4 i1_2_lut_rep_316_3_lut (.A(count[9]), .B(n13631), .C(count[8]), 
         .Z(n31460)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_316_3_lut.init = 16'hfefe;
    LUT4 i15667_2_lut_3_lut_4_lut (.A(count[9]), .B(n13631), .C(n31495), 
         .D(count[8]), .Z(n22410)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i15667_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_293_3_lut_4_lut (.A(count[9]), .B(n13631), .C(n27662), 
         .D(count[8]), .Z(n31437)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[28:39])
    defparam i1_2_lut_rep_293_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_351 (.A(n129_adj_206), .B(count[1]), .C(count[0]), 
         .Z(n31495)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_3_lut_rep_351.init = 16'h8080;
    LUT4 i1_2_lut_rep_317_4_lut (.A(n129_adj_206), .B(count[1]), .C(count[0]), 
         .D(count[8]), .Z(n31461)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_317_4_lut.init = 16'h8000;
    LUT4 i22095_3_lut_4_lut (.A(n31461), .B(n29518), .C(n31494), .D(n23), 
         .Z(n29654)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i22095_3_lut_4_lut.init = 16'hfffe;
    LUT4 i22448_3_lut_4_lut_4_lut (.A(n31482), .B(n29518), .C(n31460), 
         .D(n27662), .Z(n29398)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i22448_3_lut_4_lut_4_lut.init = 16'h1110;
    LUT4 i1_2_lut_rep_422 (.A(n1186), .B(n1174), .Z(n31566)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_422.init = 16'hbbbb;
    LUT4 i22372_2_lut_3_lut (.A(n1186), .B(n1174), .C(n27609), .Z(n29832)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i22372_2_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_426 (.A(count[5]), .B(count[4]), .Z(n31570)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_426.init = 16'h8888;
    LUT4 i2_3_lut_4_lut (.A(count[5]), .B(count[4]), .C(n29187), .D(n31599), 
         .Z(n129_adj_206)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_3_lut_4_lut.init = 16'h8000;
    IFS1P3DX latched_in_45 (.D(rc_ch2_c), .SP(n33387), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1186));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i5_2_lut_rep_429 (.A(n1174), .B(n1186), .Z(n31573)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_429.init = 16'h4444;
    LUT4 i1_2_lut_3_lut (.A(n1174), .B(n1186), .C(n31482), .Z(n29397)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut.init = 16'hf4f4;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n31412), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n31412), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n31412), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n31412), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n31412), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n31412), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n31412), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n31412), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33388), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33388), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14513), .PD(n16910), .CK(debug_c_c), 
            .Q(\register[2] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14513), .PD(n16910), .CK(debug_c_c), 
            .Q(\register[2] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14513), .PD(n16910), .CK(debug_c_c), 
            .Q(\register[2] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14513), .PD(n16910), .CK(debug_c_c), 
            .Q(\register[2] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14513), .PD(n16910), .CK(debug_c_c), 
            .Q(\register[2] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14513), .PD(n16910), .CK(debug_c_c), 
            .Q(\register[2] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14513), .PD(n16910), .CK(debug_c_c), 
            .Q(\register[2] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1186), .SP(n33387), .CK(debug_c_c), .Q(n1174));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i21_3_lut_rep_294_4_lut (.A(count[8]), .B(n31495), .C(n31494), 
         .D(n29518), .Z(n31438)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i21_3_lut_rep_294_4_lut.init = 16'h00f8;
    LUT4 i1_2_lut_3_lut_adj_291 (.A(count[8]), .B(n31495), .C(count[9]), 
         .Z(n18)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_adj_291.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_455 (.A(count[6]), .B(count[7]), .Z(n31599)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_rep_455.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_292 (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_2_lut_3_lut_adj_292.init = 16'h8080;
    LUT4 i22387_4_lut (.A(n29248), .B(n31573), .C(n31482), .D(n31566), 
         .Z(n29847)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i22387_4_lut.init = 16'h3031;
    LUT4 i3_4_lut (.A(n31460), .B(n29654), .C(n31495), .D(n27662), .Z(n29248)) /* synthesis lut_function=(!(A (B)+!A (B+!(C (D))))) */ ;
    defparam i3_4_lut.init = 16'h3222;
    FD1P3IX valid_48 (.D(n29398), .SP(n27536), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1180));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    CCU2D add_1779_17 (.A0(count[15]), .B0(n31573), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26495), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_17.INIT0 = 16'hd222;
    defparam add_1779_17.INIT1 = 16'h0000;
    defparam add_1779_17.INJECT1_0 = "NO";
    defparam add_1779_17.INJECT1_1 = "NO";
    CCU2D sub_75_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26751), 
          .S0(n1102[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_75_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_75_add_2_9.INIT1 = 16'h0000;
    defparam sub_75_add_2_9.INJECT1_0 = "NO";
    defparam sub_75_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_75_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26750), 
          .COUT(n26751), .S0(n1102[5]), .S1(n1102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_75_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_75_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_75_add_2_7.INJECT1_0 = "NO";
    defparam sub_75_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_75_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26749), 
          .COUT(n26750), .S0(n1102[3]), .S1(n1102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_75_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_75_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_75_add_2_5.INJECT1_0 = "NO";
    defparam sub_75_add_2_5.INJECT1_1 = "NO";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14513), .PD(n16910), .CK(debug_c_c), 
            .Q(\register[2] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D sub_75_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26748), 
          .COUT(n26749), .S0(n1102[1]), .S1(n1102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_75_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_75_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_75_add_2_3.INJECT1_0 = "NO";
    defparam sub_75_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_75_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26748), 
          .S1(n1102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_75_add_2_1.INIT0 = 16'hF000;
    defparam sub_75_add_2_1.INIT1 = 16'h5555;
    defparam sub_75_add_2_1.INJECT1_0 = "NO";
    defparam sub_75_add_2_1.INJECT1_1 = "NO";
    LUT4 i3_4_lut_adj_293 (.A(n33386), .B(n28999), .C(n1174), .D(n29518), 
         .Z(n16910)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_293.init = 16'h0080;
    LUT4 i3_4_lut_adj_294 (.A(n27609), .B(n1186), .C(n31512), .D(n18), 
         .Z(n28999)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_294.init = 16'h0200;
    LUT4 i15403_2_lut (.A(n1102[7]), .B(n23), .Z(n43[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15403_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(count[8]), .B(n31494), .C(count[1]), .D(n129_adj_206), 
         .Z(n23)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0222;
    LUT4 i2_4_lut_adj_295 (.A(n31438), .B(n23), .C(n31437), .D(n22410), 
         .Z(n27609)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i2_4_lut_adj_295.init = 16'heefe;
    LUT4 i2_4_lut_adj_296 (.A(n31599), .B(count[4]), .C(count[5]), .D(n4_adj_207), 
         .Z(n27662)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_296.init = 16'ha080;
    LUT4 i1_3_lut (.A(count[3]), .B(count[1]), .C(count[2]), .Z(n4_adj_207)) /* synthesis lut_function=(A+(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_3_lut.init = 16'heaea;
    LUT4 i21964_4_lut (.A(n13631), .B(count[9]), .C(n5), .D(n6), .Z(n29518)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i21964_4_lut.init = 16'heeea;
    LUT4 i1_2_lut_adj_297 (.A(count[8]), .B(count[6]), .Z(n5)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_adj_297.init = 16'heeee;
    LUT4 i2_4_lut_adj_298 (.A(count[7]), .B(count[3]), .C(n31570), .D(n27518), 
         .Z(n6)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i2_4_lut_adj_298.init = 16'hfaea;
    LUT4 i2_3_lut (.A(count[0]), .B(count[2]), .C(count[1]), .Z(n27518)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i3_4_lut_adj_299 (.A(count[12]), .B(count[13]), .C(n13702), .D(n29351), 
         .Z(n13631)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_299.init = 16'hfffe;
    LUT4 i15402_2_lut (.A(n1102[6]), .B(n23), .Z(n43[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15402_2_lut.init = 16'h8888;
    LUT4 i15401_2_lut (.A(n1102[5]), .B(n23), .Z(n43[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15401_2_lut.init = 16'h8888;
    LUT4 i15400_2_lut (.A(n1102[4]), .B(n23), .Z(n43[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15400_2_lut.init = 16'h8888;
    LUT4 i15399_2_lut (.A(n1102[3]), .B(n23), .Z(n43[3])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15399_2_lut.init = 16'h8888;
    LUT4 i15398_2_lut (.A(n1102[2]), .B(n23), .Z(n43[2])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15398_2_lut.init = 16'h8888;
    LUT4 i15397_2_lut (.A(n1102[1]), .B(n23), .Z(n43[1])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15397_2_lut.init = 16'h8888;
    LUT4 i15176_2_lut (.A(n1102[0]), .B(n23), .Z(n43[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15176_2_lut.init = 16'h8888;
    CCU2D add_1779_15 (.A0(count[13]), .B0(n31573), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n31573), .C1(GND_net), .D1(GND_net), .CIN(n26494), 
          .COUT(n26495), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_15.INIT0 = 16'hd222;
    defparam add_1779_15.INIT1 = 16'hd222;
    defparam add_1779_15.INJECT1_0 = "NO";
    defparam add_1779_15.INJECT1_1 = "NO";
    CCU2D add_1779_13 (.A0(count[11]), .B0(n31573), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n31573), .C1(GND_net), .D1(GND_net), .CIN(n26493), 
          .COUT(n26494), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_13.INIT0 = 16'hd222;
    defparam add_1779_13.INIT1 = 16'hd222;
    defparam add_1779_13.INJECT1_0 = "NO";
    defparam add_1779_13.INJECT1_1 = "NO";
    CCU2D add_1779_11 (.A0(count[9]), .B0(n31573), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n31573), .C1(GND_net), .D1(GND_net), .CIN(n26492), 
          .COUT(n26493), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_11.INIT0 = 16'hd222;
    defparam add_1779_11.INIT1 = 16'hd222;
    defparam add_1779_11.INJECT1_0 = "NO";
    defparam add_1779_11.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U5
//

module PWMReceiver_U5 (debug_c_c, n33387, \register[1] , n14514, rc_ch1_c, 
            GND_net, n29830, n33386, n1165, n27547, n29811) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n33387;
    output [7:0]\register[1] ;
    input n14514;
    input rc_ch1_c;
    input GND_net;
    output n29830;
    input n33386;
    output n1165;
    input n27547;
    output n29811;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n31577, n29366, n31496, n31579, n31580, n31578, n29287, 
        n1159, n1171, n29111, n31442, n33382, n31440, n29403, 
        n27608, n10, n31441, n31528, n31462, n28948, n7, n10_adj_204, 
        n29569, n27648, n16913;
    wire [7:0]n43;
    
    wire n5, n29404, n31529, n29110, n31527, n26503;
    wire [15:0]n116;
    
    wire n26502, n26501, n29524, n26500, n26499, n16, n26, n26498;
    wire [7:0]n1093;
    
    wire n26755, n26754, n27575, n6, n26497, n26496, n26753, n26752, 
        n6_adj_205, n4, n27503, n27546;
    
    LUT4 i3_3_lut_rep_352_4_lut (.A(count[12]), .B(n31577), .C(n29366), 
         .D(count[13]), .Z(n31496)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_3_lut_rep_352_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[0]), .B(n31579), .C(n31580), .D(n31578), 
         .Z(n29287)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1P3AX prev_in_46 (.D(n1171), .SP(n33387), .CK(debug_c_c), .Q(n1159));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i22477_3_lut_3_lut_4_lut (.A(n29111), .B(n31442), .C(n33382), 
         .D(n31440), .Z(n29403)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i22477_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i21_3_lut_rep_297_4_lut_4_lut (.A(n27608), .B(n31496), .C(count[9]), 
         .D(n10), .Z(n31441)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(C+(D))))) */ ;
    defparam i21_3_lut_rep_297_4_lut_4_lut.init = 16'h1310;
    LUT4 i22011_3_lut_rep_465 (.A(n27608), .B(n31496), .C(count[9]), .Z(n33382)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i22011_3_lut_rep_465.init = 16'hecec;
    LUT4 i1_2_lut_rep_318_4_lut (.A(n31528), .B(count[13]), .C(n29366), 
         .D(count[9]), .Z(n31462)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_318_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut (.A(n10), .B(n33382), .C(n31462), .D(n28948), 
         .Z(n7)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i1_2_lut_4_lut.init = 16'hcd00;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n31462), .C(n29287), 
         .D(n29111), .Z(n10_adj_204)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i22013_3_lut_4_lut (.A(count[8]), .B(n31462), .C(n29111), .D(n29287), 
         .Z(n29569)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i22013_3_lut_4_lut.init = 16'hfeee;
    LUT4 i1_2_lut_rep_433 (.A(count[15]), .B(count[14]), .Z(n31577)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_433.init = 16'heeee;
    LUT4 i1_2_lut_rep_296_3_lut (.A(count[15]), .B(count[14]), .C(n27648), 
         .Z(n31440)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_296_3_lut.init = 16'hfefe;
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n14514), .PD(n16913), .CK(debug_c_c), 
            .Q(\register[1] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_281 (.A(count[15]), .B(count[14]), .C(n5), 
         .D(n27648), .Z(n29404)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_281.init = 16'hfffe;
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n14514), .PD(n16913), .CK(debug_c_c), 
            .Q(\register[1] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n14514), .PD(n16913), .CK(debug_c_c), 
            .Q(\register[1] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n14514), .PD(n16913), .CK(debug_c_c), 
            .Q(\register[1] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n14514), .PD(n16913), .CK(debug_c_c), 
            .Q(\register[1] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    LUT4 i21958_2_lut_rep_384_3_lut (.A(count[15]), .B(count[14]), .C(count[12]), 
         .Z(n31528)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i21958_2_lut_rep_384_3_lut.init = 16'hfefe;
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n14514), .PD(n16913), .CK(debug_c_c), 
            .Q(\register[1] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n14514), .PD(n16913), .CK(debug_c_c), 
            .Q(\register[1] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i14717_2_lut_rep_434 (.A(count[4]), .B(count[5]), .Z(n31578)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14717_2_lut_rep_434.init = 16'h8888;
    LUT4 i2_3_lut_rep_435 (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n31579)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_rep_435.init = 16'h8080;
    LUT4 i1_2_lut_rep_385_4_lut (.A(count[2]), .B(count[3]), .C(count[1]), 
         .D(count[0]), .Z(n31529)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_385_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_436 (.A(count[6]), .B(count[7]), .Z(n31580)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_436.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[6]), .B(count[7]), .C(count[5]), .Z(n29110)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i2_2_lut_rep_383_3_lut_4_lut (.A(count[6]), .B(count[7]), .C(count[5]), 
         .D(count[4]), .Z(n31527)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_2_lut_rep_383_3_lut_4_lut.init = 16'h8000;
    IFS1P3DX latched_in_45 (.D(rc_ch1_c), .SP(n33387), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1171));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i5_2_lut (.A(n1159), .B(n1171), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_rep_298_3_lut (.A(count[9]), .B(n31496), .C(count[8]), 
         .Z(n31442)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_298_3_lut.init = 16'hfefe;
    CCU2D add_1775_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26503), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_17.INIT0 = 16'hd222;
    defparam add_1775_17.INIT1 = 16'h0000;
    defparam add_1775_17.INJECT1_0 = "NO";
    defparam add_1775_17.INJECT1_1 = "NO";
    CCU2D add_1775_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26502), 
          .COUT(n26503), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_15.INIT0 = 16'hd222;
    defparam add_1775_15.INIT1 = 16'hd222;
    defparam add_1775_15.INJECT1_0 = "NO";
    defparam add_1775_15.INJECT1_1 = "NO";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    CCU2D add_1775_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26501), 
          .COUT(n26502), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_13.INIT0 = 16'hd222;
    defparam add_1775_13.INIT1 = 16'hd222;
    defparam add_1775_13.INJECT1_0 = "NO";
    defparam add_1775_13.INJECT1_1 = "NO";
    LUT4 i22370_4_lut (.A(n31441), .B(n29524), .C(n28948), .D(n10_adj_204), 
         .Z(n29830)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i22370_4_lut.init = 16'h3323;
    CCU2D add_1775_11 (.A0(count[9]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26500), 
          .COUT(n26501), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_11.INIT0 = 16'hd222;
    defparam add_1775_11.INIT1 = 16'hd222;
    defparam add_1775_11.INJECT1_0 = "NO";
    defparam add_1775_11.INJECT1_1 = "NO";
    CCU2D add_1775_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26499), 
          .COUT(n26500), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_9.INIT0 = 16'hd222;
    defparam add_1775_9.INIT1 = 16'hd222;
    defparam add_1775_9.INJECT1_0 = "NO";
    defparam add_1775_9.INJECT1_1 = "NO";
    LUT4 i8_4_lut (.A(n31528), .B(n16), .C(count[13]), .D(count[11]), 
         .Z(n16913)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i8_4_lut.init = 16'h0004;
    LUT4 i7_4_lut (.A(count[10]), .B(n33386), .C(n26), .D(n29524), .Z(n16)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i7_4_lut.init = 16'h0040;
    CCU2D add_1775_7 (.A0(count[5]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26498), 
          .COUT(n26499), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_7.INIT0 = 16'hd222;
    defparam add_1775_7.INIT1 = 16'hd222;
    defparam add_1775_7.INJECT1_0 = "NO";
    defparam add_1775_7.INJECT1_1 = "NO";
    LUT4 i33_3_lut (.A(n10), .B(n27608), .C(count[9]), .Z(n26)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i33_3_lut.init = 16'h3a3a;
    LUT4 i15396_2_lut (.A(n1093[7]), .B(n28948), .Z(n43[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15396_2_lut.init = 16'h2222;
    CCU2D sub_74_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26755), 
          .S0(n1093[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_74_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_74_add_2_9.INIT1 = 16'h0000;
    defparam sub_74_add_2_9.INJECT1_0 = "NO";
    defparam sub_74_add_2_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(n31462), .B(count[8]), .C(n31579), .D(n31527), 
         .Z(n28948)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfbbb;
    LUT4 i3_4_lut (.A(count[4]), .B(n31529), .C(count[8]), .D(n29110), 
         .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut.init = 16'h8000;
    CCU2D sub_74_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26754), 
          .COUT(n26755), .S0(n1093[5]), .S1(n1093[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_74_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_74_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_74_add_2_7.INJECT1_0 = "NO";
    defparam sub_74_add_2_7.INJECT1_1 = "NO";
    LUT4 i3_4_lut_adj_282 (.A(n27575), .B(n6), .C(count[8]), .D(n31578), 
         .Z(n27608)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_282.init = 16'hfefc;
    LUT4 i3_4_lut_adj_283 (.A(count[0]), .B(count[1]), .C(count[3]), .D(count[2]), 
         .Z(n27575)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_283.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[6]), .B(count[7]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    CCU2D add_1775_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26497), 
          .COUT(n26498), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_5.INIT0 = 16'hd222;
    defparam add_1775_5.INIT1 = 16'hd222;
    defparam add_1775_5.INJECT1_0 = "NO";
    defparam add_1775_5.INJECT1_1 = "NO";
    CCU2D add_1775_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n26496), 
          .COUT(n26497), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_3.INIT0 = 16'hd222;
    defparam add_1775_3.INIT1 = 16'hd222;
    defparam add_1775_3.INJECT1_0 = "NO";
    defparam add_1775_3.INJECT1_1 = "NO";
    CCU2D sub_74_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26753), 
          .COUT(n26754), .S0(n1093[3]), .S1(n1093[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_74_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_74_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_74_add_2_5.INJECT1_0 = "NO";
    defparam sub_74_add_2_5.INJECT1_1 = "NO";
    CCU2D add_1775_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n29404), .B1(n1171), .C1(count[0]), .D1(n1159), .COUT(n26496), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_1.INIT0 = 16'hF000;
    defparam add_1775_1.INIT1 = 16'ha565;
    defparam add_1775_1.INJECT1_0 = "NO";
    defparam add_1775_1.INJECT1_1 = "NO";
    CCU2D sub_74_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n26752), 
          .COUT(n26753), .S0(n1093[1]), .S1(n1093[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_74_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_74_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_74_add_2_3.INJECT1_0 = "NO";
    defparam sub_74_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_74_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n26752), 
          .S1(n1093[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_74_add_2_1.INIT0 = 16'hF000;
    defparam sub_74_add_2_1.INIT1 = 16'h5555;
    defparam sub_74_add_2_1.INJECT1_0 = "NO";
    defparam sub_74_add_2_1.INJECT1_1 = "NO";
    LUT4 i21970_2_lut (.A(n1159), .B(n1171), .Z(n29524)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i21970_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut (.A(count[11]), .B(count[10]), .Z(n29366)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_284 (.A(count[4]), .B(n29110), .C(count[3]), .D(n6_adj_205), 
         .Z(n29111)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_284.init = 16'hccc8;
    LUT4 i3301_2_lut (.A(count[1]), .B(count[2]), .Z(n6_adj_205)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3301_2_lut.init = 16'h8888;
    LUT4 i15395_2_lut (.A(n1093[6]), .B(n28948), .Z(n43[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15395_2_lut.init = 16'h2222;
    LUT4 i15394_2_lut (.A(n1093[5]), .B(n28948), .Z(n43[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15394_2_lut.init = 16'h2222;
    LUT4 i15393_2_lut (.A(n1093[4]), .B(n28948), .Z(n43[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15393_2_lut.init = 16'h2222;
    LUT4 i15392_2_lut (.A(n1093[3]), .B(n28948), .Z(n43[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15392_2_lut.init = 16'h2222;
    FD1P3AX valid_48 (.D(n29403), .SP(n27547), .CK(debug_c_c), .Q(n1165));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n14514), .PD(n16913), .CK(debug_c_c), 
            .Q(\register[1] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n29366), .D(n4), 
         .Z(n27648)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_4_lut_adj_285 (.A(n31580), .B(count[9]), .C(n27503), .D(count[8]), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_285.init = 16'heccc;
    LUT4 i2_4_lut_adj_286 (.A(count[5]), .B(count[4]), .C(n6_adj_205), 
         .D(count[3]), .Z(n27503)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_286.init = 16'hfeee;
    LUT4 i15391_2_lut (.A(n1093[2]), .B(n28948), .Z(n43[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15391_2_lut.init = 16'h2222;
    LUT4 i15390_2_lut (.A(n1093[1]), .B(n28948), .Z(n43[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15390_2_lut.init = 16'h2222;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n33387), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    LUT4 i22351_4_lut (.A(n31577), .B(n5), .C(n27648), .D(n27546), .Z(n29811)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i22351_4_lut.init = 16'h3233;
    LUT4 i1_4_lut_adj_287 (.A(n33382), .B(n29524), .C(n7), .D(n29569), 
         .Z(n27546)) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_287.init = 16'hdccc;
    LUT4 i15173_2_lut (.A(n1093[0]), .B(n28948), .Z(n43[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15173_2_lut.init = 16'h2222;
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n33387), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module SabertoothSerialPeripheral
//

module SabertoothSerialPeripheral (\read_size[0] , debug_c_c, n9379, n13908, 
            n31512, \databus[0] , \select[2] , read_value, n9542, 
            rw, n64, n31601, \register[0][7] , n31582, \reset_count[14] , 
            n22484, n11236, \databus[7] , \databus[6] , \databus[5] , 
            \databus[4] , \databus[3] , \databus[2] , \databus[1] , 
            \register_addr[0] , n31413, GND_net, n1156, n31537, \reset_count[8] , 
            \reset_count[7] , n29332, state, n29170, n31596, n31556, 
            n31576, n9, n33385, n31443, n31590, n35, n4181, \register_addr[5] , 
            n31464, n13917, \reset_count[11] , n21503, n27250, n29264, 
            n14783, n31530, n9297, n31463, n11073, n8507, n29786, 
            select_clk, n2967, n107) /* synthesis syn_module_defined=1 */ ;
    output \read_size[0] ;
    input debug_c_c;
    input n9379;
    input n13908;
    input n31512;
    input \databus[0] ;
    input \select[2] ;
    output [7:0]read_value;
    input n9542;
    input rw;
    output n64;
    input n31601;
    output \register[0][7] ;
    output n31582;
    input \reset_count[14] ;
    input n22484;
    input n11236;
    input \databus[7] ;
    input \databus[6] ;
    input \databus[5] ;
    input \databus[4] ;
    input \databus[3] ;
    input \databus[2] ;
    input \databus[1] ;
    input \register_addr[0] ;
    input n31413;
    input GND_net;
    output n1156;
    input n31537;
    input \reset_count[8] ;
    input \reset_count[7] ;
    output n29332;
    output [3:0]state;
    input n29170;
    input n31596;
    input n31556;
    input n31576;
    output n9;
    input n33385;
    input n31443;
    input n31590;
    input n35;
    output n4181;
    input \register_addr[5] ;
    input n31464;
    output n13917;
    input \reset_count[11] ;
    input n21503;
    input n27250;
    output n29264;
    input n14783;
    input n31530;
    output n9297;
    input n31463;
    output n11073;
    output n8507;
    output n29786;
    output select_clk;
    input n2967;
    input n107;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n14967;
    wire [7:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    
    wire prev_select;
    wire [7:0]n28;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    
    wire n29474, n9449;
    wire [31:0]n63;
    
    wire n31534, n27245, n9446;
    wire [7:0]n6205;
    
    FD1P3AX read_size__i1 (.D(n9379), .SP(n14967), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3JX register_0__i1 (.D(\databus[0] ), .SP(n13908), .PD(n31512), 
            .CK(debug_c_c), .Q(\register[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i1.GSR = "ENABLED";
    FD1S3AX prev_select_138 (.D(\select[2] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam prev_select_138.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n28[0]), .SP(n14967), .CD(n9542), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i16_2_lut (.A(\select[2] ), .B(rw), .Z(n64)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(97[19:32])
    defparam i16_2_lut.init = 16'h8888;
    LUT4 i15388_4_lut_4_lut (.A(\register[1] [7]), .B(n31601), .C(n29474), 
         .D(n9449), .Z(n63[6])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(89[23:51])
    defparam i15388_4_lut_4_lut.init = 16'hffde;
    LUT4 i1_4_lut_4_lut (.A(\register[1] [7]), .B(n31601), .C(\register[1] [1]), 
         .D(n31534), .Z(n9449)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(89[23:51])
    defparam i1_4_lut_4_lut.init = 16'h2000;
    LUT4 i1_4_lut_4_lut_adj_280 (.A(\register[0][7] ), .B(n31601), .C(\register[0] [1]), 
         .D(n27245), .Z(n9446)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(88[22:50])
    defparam i1_4_lut_4_lut_adj_280.init = 16'h2000;
    LUT4 i1_2_lut_rep_438 (.A(\select[2] ), .B(prev_select), .Z(n31582)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(110[8:29])
    defparam i1_2_lut_rep_438.init = 16'h2222;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(\select[2] ), .B(prev_select), .C(\reset_count[14] ), 
         .D(n22484), .Z(n14967)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(110[8:29])
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'h2000;
    FD1P3IX register_0__i16 (.D(\databus[7] ), .SP(n11236), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i16.GSR = "ENABLED";
    FD1P3JX register_0__i15 (.D(\databus[6] ), .SP(n11236), .PD(n31512), 
            .CK(debug_c_c), .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i15.GSR = "ENABLED";
    FD1P3JX register_0__i14 (.D(\databus[5] ), .SP(n11236), .PD(n31512), 
            .CK(debug_c_c), .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i14.GSR = "ENABLED";
    FD1P3JX register_0__i13 (.D(\databus[4] ), .SP(n11236), .PD(n31512), 
            .CK(debug_c_c), .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i13.GSR = "ENABLED";
    FD1P3JX register_0__i12 (.D(\databus[3] ), .SP(n11236), .PD(n31512), 
            .CK(debug_c_c), .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i12.GSR = "ENABLED";
    FD1P3JX register_0__i11 (.D(\databus[2] ), .SP(n11236), .PD(n31512), 
            .CK(debug_c_c), .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i11.GSR = "ENABLED";
    FD1P3JX register_0__i10 (.D(\databus[1] ), .SP(n11236), .PD(n31512), 
            .CK(debug_c_c), .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i10.GSR = "ENABLED";
    FD1P3JX register_0__i9 (.D(\databus[0] ), .SP(n11236), .PD(n31512), 
            .CK(debug_c_c), .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i9.GSR = "ENABLED";
    FD1P3IX register_0__i8 (.D(\databus[7] ), .SP(n13908), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[0][7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i8.GSR = "ENABLED";
    FD1P3JX register_0__i7 (.D(\databus[6] ), .SP(n13908), .PD(n31512), 
            .CK(debug_c_c), .Q(\register[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i7.GSR = "ENABLED";
    FD1P3JX register_0__i6 (.D(\databus[5] ), .SP(n13908), .PD(n31512), 
            .CK(debug_c_c), .Q(\register[0] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i6.GSR = "ENABLED";
    FD1P3JX register_0__i5 (.D(\databus[4] ), .SP(n13908), .PD(n31512), 
            .CK(debug_c_c), .Q(\register[0] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i5.GSR = "ENABLED";
    FD1P3JX register_0__i4 (.D(\databus[3] ), .SP(n13908), .PD(n31512), 
            .CK(debug_c_c), .Q(\register[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i4.GSR = "ENABLED";
    FD1P3JX register_0__i3 (.D(\databus[2] ), .SP(n13908), .PD(n31512), 
            .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i3.GSR = "ENABLED";
    FD1P3JX register_0__i2 (.D(\databus[1] ), .SP(n13908), .PD(n31512), 
            .CK(debug_c_c), .Q(\register[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i2.GSR = "ENABLED";
    LUT4 mux_1916_Mux_7_i1_3_lut (.A(\register[0][7] ), .B(\register[1] [7]), 
         .C(\register_addr[0] ), .Z(n6205[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1916_Mux_7_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1916_Mux_6_i1_3_lut (.A(\register[0] [6]), .B(\register[1] [6]), 
         .C(\register_addr[0] ), .Z(n6205[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1916_Mux_6_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1916_Mux_5_i1_3_lut (.A(\register[0] [5]), .B(\register[1] [5]), 
         .C(\register_addr[0] ), .Z(n6205[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1916_Mux_5_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1916_Mux_4_i1_3_lut (.A(\register[0] [4]), .B(\register[1] [4]), 
         .C(\register_addr[0] ), .Z(n6205[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1916_Mux_4_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1916_Mux_3_i1_3_lut (.A(\register[0] [3]), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n6205[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1916_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1916_Mux_2_i1_3_lut (.A(\register[0] [2]), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n6205[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1916_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1916_Mux_1_i1_3_lut (.A(\register[0] [1]), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n6205[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1916_Mux_1_i1_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i7 (.D(n6205[7]), .SP(n14967), .CD(n9542), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6205[6]), .SP(n14967), .CD(n9542), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n6205[5]), .SP(n14967), .CD(n9542), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6205[4]), .SP(n14967), .CD(n9542), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6205[3]), .SP(n14967), .CD(n9542), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n6205[2]), .SP(n14967), .CD(n9542), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n6205[1]), .SP(n14967), .CD(n9542), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 mux_1916_Mux_0_i1_3_lut (.A(\register[0] [0]), .B(\register[1] [0]), 
         .C(\register_addr[0] ), .Z(n28[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1916_Mux_0_i1_3_lut.init = 16'hcaca;
    SabertoothSerial sserial (.debug_c_c(debug_c_c), .n31413(n31413), .GND_net(GND_net), 
            .\register[0][5] (\register[0] [5]), .n31601(n31601), .\register[0][6] (\register[0] [6]), 
            .\register[1][6] (\register[1] [6]), .n31534(n31534), .\register[1][7] (\register[1] [7]), 
            .\register[1][1] (\register[1] [1]), .\register[1][3] (\register[1] [3]), 
            .\register[1][5] (\register[1] [5]), .\register[1][4] (\register[1] [4]), 
            .\register[0][3] (\register[0] [3]), .\register[0][4] (\register[0] [4]), 
            .n1156(n1156), .n29474(n29474), .n89(n63[6]), .\register[0][7] (\register[0][7] ), 
            .n9446(n9446), .\register[1][2] (\register[1] [2]), .\register[0][2] (\register[0] [2]), 
            .n27245(n27245), .n31537(n31537), .n9449(n9449), .\register[0][1] (\register[0] [1]), 
            .\reset_count[8] (\reset_count[8] ), .\reset_count[7] (\reset_count[7] ), 
            .n29332(n29332), .state({state}), .n31512(n31512), .n29170(n29170), 
            .n31596(n31596), .n31556(n31556), .n31576(n31576), .n9(n9), 
            .n33385(n33385), .n31443(n31443), .n31590(n31590), .n35(n35), 
            .n4181(n4181), .rw(rw), .\register_addr[5] (\register_addr[5] ), 
            .n31464(n31464), .n13917(n13917), .\reset_count[11] (\reset_count[11] ), 
            .n21503(n21503), .n27250(n27250), .n29264(n29264), .n14783(n14783), 
            .n31530(n31530), .n9297(n9297), .n31463(n31463), .n11073(n11073), 
            .n22484(n22484), .\reset_count[14] (\reset_count[14] ), .n8507(n8507), 
            .n29786(n29786), .select_clk(select_clk), .n2967(n2967), .n107(n107)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(142[19] 147[34])
    
endmodule
//
// Verilog Description of module SabertoothSerial
//

module SabertoothSerial (debug_c_c, n31413, GND_net, \register[0][5] , 
            n31601, \register[0][6] , \register[1][6] , n31534, \register[1][7] , 
            \register[1][1] , \register[1][3] , \register[1][5] , \register[1][4] , 
            \register[0][3] , \register[0][4] , n1156, n29474, n89, 
            \register[0][7] , n9446, \register[1][2] , \register[0][2] , 
            n27245, n31537, n9449, \register[0][1] , \reset_count[8] , 
            \reset_count[7] , n29332, state, n31512, n29170, n31596, 
            n31556, n31576, n9, n33385, n31443, n31590, n35, n4181, 
            rw, \register_addr[5] , n31464, n13917, \reset_count[11] , 
            n21503, n27250, n29264, n14783, n31530, n9297, n31463, 
            n11073, n22484, \reset_count[14] , n8507, n29786, select_clk, 
            n2967, n107) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n31413;
    input GND_net;
    input \register[0][5] ;
    input n31601;
    input \register[0][6] ;
    input \register[1][6] ;
    output n31534;
    input \register[1][7] ;
    input \register[1][1] ;
    input \register[1][3] ;
    input \register[1][5] ;
    input \register[1][4] ;
    input \register[0][3] ;
    input \register[0][4] ;
    output n1156;
    output n29474;
    input n89;
    input \register[0][7] ;
    input n9446;
    input \register[1][2] ;
    input \register[0][2] ;
    output n27245;
    input n31537;
    input n9449;
    input \register[0][1] ;
    input \reset_count[8] ;
    input \reset_count[7] ;
    output n29332;
    output [3:0]state;
    input n31512;
    input n29170;
    input n31596;
    input n31556;
    input n31576;
    output n9;
    input n33385;
    input n31443;
    input n31590;
    input n35;
    output n4181;
    input rw;
    input \register_addr[5] ;
    input n31464;
    output n13917;
    input \reset_count[11] ;
    input n21503;
    input n27250;
    output n29264;
    input n14783;
    input n31530;
    output n9297;
    input n31463;
    output n11073;
    input n22484;
    input \reset_count[14] ;
    output n8507;
    output n29786;
    output select_clk;
    input n2967;
    input n107;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [3:0]state_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(17[12:17])
    wire [3:0]n7809;
    wire [3:0]n16;
    
    wire n1, n31505, n10325;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(16[12:19])
    
    wire n14037, n31405, n29224, n20, n31587, n31472, n31589, 
        n31475, n12743, n31536, n31538, n12741, n28954, n6, n7, 
        n28311, n8;
    wire [7:0]n5505;
    wire [7:0]n5514;
    
    wire n12_adj_199;
    wire [31:0]n63;
    
    wire n6_adj_200, n11382, n11964, n12016, n12134, n24, n31503;
    
    FD1P3IX state__i1 (.D(n7809[1]), .SP(n31413), .CD(GND_net), .CK(debug_c_c), 
            .Q(state_c[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam state__i1.GSR = "ENABLED";
    FD1S3IX state__i0 (.D(n16[0]), .CK(debug_c_c), .CD(GND_net), .Q(state_c[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam state__i0.GSR = "ENABLED";
    LUT4 i3948_1_lut (.A(state_c[0]), .Z(n1)) /* synthesis lut_function=(!(A)) */ ;
    defparam i3948_1_lut.init = 16'h5555;
    LUT4 i15445_3_lut_4_lut (.A(\register[0][5] ), .B(n31505), .C(n31601), 
         .D(\register[0][6] ), .Z(n10325)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i15445_3_lut_4_lut.init = 16'hf8f0;
    FD1P3AX tx_data_i0_i0 (.D(n31405), .SP(n14037), .CK(debug_c_c), .Q(tx_data[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_390 (.A(\register[1][6] ), .B(n29224), .Z(n31534)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_390.init = 16'h8888;
    LUT4 i1_3_lut_4_lut (.A(\register[1][6] ), .B(n29224), .C(\register[1][7] ), 
         .D(\register[1][1] ), .Z(n20)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h80ff;
    LUT4 i5806_2_lut_rep_328_3_lut_4_lut (.A(\register[1][3] ), .B(n31587), 
         .C(\register[1][5] ), .D(\register[1][4] ), .Z(n31472)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5806_2_lut_rep_328_3_lut_4_lut.init = 16'h8000;
    LUT4 i5958_2_lut_rep_331_3_lut_4_lut (.A(\register[0][3] ), .B(n31589), 
         .C(\register[0][5] ), .D(\register[0][4] ), .Z(n31475)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5958_2_lut_rep_331_3_lut_4_lut.init = 16'h8000;
    LUT4 i5974_2_lut_3_lut_4_lut (.A(\register[0][3] ), .B(n31589), .C(\register[0][5] ), 
         .D(\register[0][4] ), .Z(n12743)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i5974_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1P3IX send_31 (.D(n1), .SP(n31413), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1156));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam send_31.GSR = "ENABLED";
    LUT4 i4377_2_lut (.A(state_c[0]), .B(state_c[1]), .Z(n7809[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(34[6] 57[13])
    defparam i4377_2_lut.init = 16'h6666;
    LUT4 i21922_2_lut_3_lut_4_lut (.A(\register[1][4] ), .B(n31536), .C(\register[1][6] ), 
         .D(\register[1][5] ), .Z(n29474)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i21922_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i5972_2_lut_3_lut_4_lut (.A(\register[0][4] ), .B(n31538), .C(\register[0][6] ), 
         .D(\register[0][5] ), .Z(n12741)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i5972_2_lut_3_lut_4_lut.init = 16'h78f0;
    PFUMX i30 (.BLUT(n28954), .ALUT(n6), .C0(n7), .Z(n28311));
    LUT4 i1_4_lut (.A(n31601), .B(\register[1][7] ), .C(n29474), .D(n8), 
         .Z(n28954)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_4_lut.init = 16'hffbf;
    LUT4 i1_2_lut (.A(\register[1][1] ), .B(n29224), .Z(n8)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    PFUMX mux_1849_i7 (.BLUT(n89), .ALUT(n5505[6]), .C0(n7), .Z(n5514[6]));
    LUT4 i6_4_lut (.A(n31475), .B(n12_adj_199), .C(\register[0][7] ), 
         .D(state_c[1]), .Z(n6)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i6_4_lut.init = 16'h0080;
    PFUMX mux_1849_i2 (.BLUT(n63[1]), .ALUT(n5505[1]), .C0(n7), .Z(n5514[1]));
    LUT4 i5_4_lut (.A(\register[0][6] ), .B(state_c[0]), .C(n9446), .D(n31601), 
         .Z(n12_adj_199)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i5_4_lut.init = 16'h0002;
    PFUMX mux_1849_i3 (.BLUT(n63[2]), .ALUT(n5505[2]), .C0(n7), .Z(n5514[2]));
    LUT4 equal_16_i5_2_lut (.A(state_c[0]), .B(state_c[1]), .Z(n7)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(46[7:11])
    defparam equal_16_i5_2_lut.init = 16'hbbbb;
    LUT4 i3_4_lut (.A(\register[1][4] ), .B(\register[1][3] ), .C(\register[1][5] ), 
         .D(\register[1][2] ), .Z(n29224)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    PFUMX mux_1849_i4 (.BLUT(n63[3]), .ALUT(n5505[3]), .C0(n7), .Z(n5514[3]));
    LUT4 i4_4_lut (.A(\register[0][4] ), .B(\register[0][2] ), .C(\register[0][3] ), 
         .D(n6_adj_200), .Z(n27245)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i4_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_adj_278 (.A(\register[0][5] ), .B(\register[0][6] ), .Z(n6_adj_200)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_278.init = 16'h8888;
    PFUMX mux_1849_i5 (.BLUT(n63[4]), .ALUT(n5505[4]), .C0(n7), .Z(n5514[4]));
    PFUMX mux_1849_i6 (.BLUT(n63[5]), .ALUT(n5505[5]), .C0(n7), .Z(n5514[5]));
    LUT4 i15047_4_lut (.A(n31537), .B(n11382), .C(n9446), .D(n10325), 
         .Z(n5505[6])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C+(D))))) */ ;
    defparam i15047_4_lut.init = 16'h3132;
    LUT4 i4392_2_lut (.A(state_c[0]), .B(state_c[1]), .Z(n11382)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i4392_2_lut.init = 16'heeee;
    LUT4 i15383_4_lut (.A(\register[1][2] ), .B(n9449), .C(n31601), .D(\register[1][1] ), 
         .Z(n63[1])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15383_4_lut.init = 16'hcdce;
    LUT4 i15039_4_lut (.A(n11964), .B(n11382), .C(n9446), .D(n31601), 
         .Z(n5505[1])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i15039_4_lut.init = 16'h3032;
    LUT4 i5199_2_lut (.A(\register[0][2] ), .B(\register[0][1] ), .Z(n11964)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5199_2_lut.init = 16'h6666;
    LUT4 i15384_4_lut (.A(\register[1][3] ), .B(n9449), .C(n31601), .D(n31587), 
         .Z(n63[2])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15384_4_lut.init = 16'hcdce;
    LUT4 i15040_4_lut (.A(n12016), .B(n11382), .C(n9446), .D(n31601), 
         .Z(n5505[2])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i15040_4_lut.init = 16'h3032;
    LUT4 i15385_4_lut (.A(\register[1][4] ), .B(n9449), .C(n31601), .D(n31536), 
         .Z(n63[3])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15385_4_lut.init = 16'hcdce;
    LUT4 i15041_4_lut (.A(n12134), .B(n11382), .C(n9446), .D(n31601), 
         .Z(n5505[3])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i15041_4_lut.init = 16'h3032;
    LUT4 n20_bdd_4_lut (.A(n20), .B(n24), .C(n7), .D(n31601), .Z(n31405)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n20_bdd_4_lut.init = 16'h00ca;
    LUT4 i15386_4_lut (.A(\register[1][5] ), .B(n9449), .C(n31601), .D(n31503), 
         .Z(n63[4])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15386_4_lut.init = 16'hcdce;
    LUT4 i15042_4_lut (.A(n12743), .B(n11382), .C(n9446), .D(n31601), 
         .Z(n5505[4])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i15042_4_lut.init = 16'h3032;
    LUT4 i15387_4_lut (.A(\register[1][6] ), .B(n9449), .C(n31601), .D(n31472), 
         .Z(n63[5])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15387_4_lut.init = 16'hcdce;
    LUT4 i4423_2_lut_rep_443 (.A(\register[1][2] ), .B(\register[1][1] ), 
         .Z(n31587)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4423_2_lut_rep_443.init = 16'h8888;
    LUT4 i5801_2_lut_rep_359_3_lut_4_lut (.A(\register[1][2] ), .B(\register[1][1] ), 
         .C(\register[1][4] ), .D(\register[1][3] ), .Z(n31503)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5801_2_lut_rep_359_3_lut_4_lut.init = 16'h8000;
    LUT4 i15044_4_lut (.A(n12741), .B(n11382), .C(n9446), .D(n31601), 
         .Z(n5505[5])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i15044_4_lut.init = 16'h3032;
    LUT4 i4435_2_lut_rep_392_3_lut (.A(\register[1][2] ), .B(\register[1][1] ), 
         .C(\register[1][3] ), .Z(n31536)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i4435_2_lut_rep_392_3_lut.init = 16'h8080;
    LUT4 i5237_2_lut_rep_445 (.A(\register[0][2] ), .B(\register[0][1] ), 
         .Z(n31589)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5237_2_lut_rep_445.init = 16'h8888;
    LUT4 i5239_2_lut_rep_394_3_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][3] ), .Z(n31538)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5239_2_lut_rep_394_3_lut.init = 16'h8080;
    LUT4 i5251_2_lut_3_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][3] ), .Z(n12016)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i5251_2_lut_3_lut.init = 16'h7878;
    LUT4 i5956_2_lut_rep_361_3_lut_4_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][4] ), .D(\register[0][3] ), .Z(n31505)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5956_2_lut_rep_361_3_lut_4_lut.init = 16'h8000;
    LUT4 i5369_2_lut_3_lut_4_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][4] ), .D(\register[0][3] ), .Z(n12134)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i5369_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1P3AX tx_data_i0_i1 (.D(n5514[1]), .SP(n14037), .CK(debug_c_c), 
            .Q(tx_data[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i2 (.D(n5514[2]), .SP(n14037), .CK(debug_c_c), 
            .Q(tx_data[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n5514[3]), .SP(n14037), .CK(debug_c_c), 
            .Q(tx_data[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i4 (.D(n5514[4]), .SP(n14037), .CK(debug_c_c), 
            .Q(tx_data[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i5 (.D(n5514[5]), .SP(n14037), .CK(debug_c_c), 
            .Q(tx_data[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i6 (.D(n5514[6]), .SP(n14037), .CK(debug_c_c), 
            .Q(tx_data[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i7 (.D(n28311), .SP(n14037), .CK(debug_c_c), .Q(tx_data[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_279 (.A(n11382), .B(\register[0][1] ), .C(n27245), 
         .D(\register[0][7] ), .Z(n24)) /* synthesis lut_function=(!(A+!((C (D))+!B))) */ ;
    defparam i1_4_lut_adj_279.init = 16'h5111;
    \UARTTransmitter(baud_div=1250)  sender (.\reset_count[8] (\reset_count[8] ), 
            .\reset_count[7] (\reset_count[7] ), .n29332(n29332), .state({state}), 
            .n31512(n31512), .n29170(n29170), .n31596(n31596), .n31556(n31556), 
            .n31576(n31576), .n9(n9), .n33385(n33385), .n31443(n31443), 
            .n31590(n31590), .n35(n35), .n4181(n4181), .rw(rw), .\register_addr[5] (\register_addr[5] ), 
            .n31464(n31464), .n13917(n13917), .\reset_count[11] (\reset_count[11] ), 
            .n21503(n21503), .n27250(n27250), .n29264(n29264), .tx_data({tx_data}), 
            .n1156(n1156), .n14783(n14783), .n31530(n31530), .n9297(n9297), 
            .n31463(n31463), .n11073(n11073), .n22484(n22484), .\reset_count[14] (\reset_count[14] ), 
            .GND_net(GND_net), .debug_c_c(debug_c_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(63[26] 67[47])
    \ClockDividerP(factor=12000)  baud_gen (.GND_net(GND_net), .n8507(n8507), 
            .n29786(n29786), .n31512(n31512), .select_clk(select_clk), 
            .\state[0] (state_c[0]), .n14037(n14037), .n12(n16[0]), .debug_c_c(debug_c_c), 
            .n2967(n2967), .n107(n107)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(21[25] 23[48])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=1250) 
//

module \UARTTransmitter(baud_div=1250)  (\reset_count[8] , \reset_count[7] , 
            n29332, state, n31512, n29170, n31596, n31556, n31576, 
            n9, n33385, n31443, n31590, n35, n4181, rw, \register_addr[5] , 
            n31464, n13917, \reset_count[11] , n21503, n27250, n29264, 
            tx_data, n1156, n14783, n31530, n9297, n31463, n11073, 
            n22484, \reset_count[14] , GND_net, debug_c_c) /* synthesis syn_module_defined=1 */ ;
    input \reset_count[8] ;
    input \reset_count[7] ;
    output n29332;
    output [3:0]state;
    input n31512;
    input n29170;
    input n31596;
    input n31556;
    input n31576;
    output n9;
    input n33385;
    input n31443;
    input n31590;
    input n35;
    output n4181;
    input rw;
    input \register_addr[5] ;
    input n31464;
    output n13917;
    input \reset_count[11] ;
    input n21503;
    input n27250;
    output n29264;
    input [7:0]tx_data;
    input n1156;
    input n14783;
    input n31530;
    output n9297;
    input n31463;
    output n11073;
    input n22484;
    input \reset_count[14] ;
    input GND_net;
    input debug_c_c;
    
    wire bclk /* synthesis SET_AS_NETWORK=\motor_serial/sserial/sender/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n30719, n2781, n28471, n17, n30718, n30717;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n9453, n7, n10, n104, n29771, n29772, n2, n29773, n29191, 
        n29192, n10_adj_198;
    
    LUT4 i1_2_lut (.A(\reset_count[8] ), .B(\reset_count[7] ), .Z(n29332)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1S3IX state__i0 (.D(n30719), .CK(bclk), .CD(n31512), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n31512), .B(state[3]), .C(state[2]), .D(n2781), 
         .Z(n28471)) /* synthesis lut_function=(!(A+(B (C)+!B !(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i1_4_lut.init = 16'h1404;
    LUT4 i3_2_lut_4_lut (.A(n29170), .B(n31596), .C(n31556), .D(n31576), 
         .Z(n9)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i3_2_lut_4_lut.init = 16'h0200;
    LUT4 i27_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), .D(state[3]), 
         .Z(n17)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B !(C+(D))))) */ ;
    defparam i27_4_lut_4_lut.init = 16'h15fe;
    LUT4 i2_3_lut_4_lut (.A(n33385), .B(n31443), .C(n31590), .D(n35), 
         .Z(n4181)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0400;
    LUT4 i2_3_lut_4_lut_adj_274 (.A(rw), .B(n31443), .C(\register_addr[5] ), 
         .D(n31464), .Z(n13917)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i2_3_lut_4_lut_adj_274.init = 16'h0004;
    PFUMX i22646 (.BLUT(n30718), .ALUT(n30717), .C0(state[2]), .Z(n30719));
    LUT4 i1_4_lut_adj_275 (.A(\reset_count[11] ), .B(n21503), .C(\reset_count[8] ), 
         .D(n27250), .Z(n29264)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_275.init = 16'h8880;
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n9453), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    PFUMX Mux_22_i15 (.BLUT(n7), .ALUT(n10), .C0(state[3]), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;
    LUT4 state_1__bdd_2_lut (.A(state[3]), .B(state[0]), .Z(n30717)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_1__bdd_2_lut.init = 16'h1111;
    LUT4 state_1__bdd_4_lut (.A(state[1]), .B(state[3]), .C(state[0]), 
         .D(n1156), .Z(n30718)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(B (C)+!B (C+!(D)))) */ ;
    defparam state_1__bdd_4_lut.init = 16'h8f0e;
    LUT4 i22211_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n29771)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22211_3_lut.init = 16'hcaca;
    LUT4 i22212_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n29772)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22212_3_lut.init = 16'hcaca;
    LUT4 Mux_22_i7_4_lut (.A(n2), .B(n29773), .C(state[2]), .D(state[1]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i15422_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i15422_4_lut.init = 16'hfcee;
    FD1P3AX state__i3 (.D(n28471), .SP(n14783), .CK(bclk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut (.A(n31512), .B(state[2]), .C(state[3]), .D(n2781), 
         .Z(n29191)) /* synthesis lut_function=(!(A+(B (C+(D))+!B !(D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h1104;
    LUT4 i4_4_lut (.A(n31443), .B(n31530), .C(n31590), .D(rw), .Z(n9297)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i4_4_lut.init = 16'h0008;
    FD1P3AX state__i2 (.D(n29191), .SP(n14783), .CK(bclk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    FD1P3AX state__i1 (.D(n29192), .SP(n14783), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    LUT4 i1_3_lut (.A(state[1]), .B(n31463), .C(state[0]), .Z(n29192)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4848;
    FD1P3JX tx_35 (.D(n104), .SP(n17), .PD(n31512), .CK(bclk), .Q(n11073)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    PFUMX i22213 (.BLUT(n29771), .ALUT(n29772), .C0(state[1]), .Z(n29773));
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n9453), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n9453), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n9453), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n9453), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n9453), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n9453), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n9453), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_276 (.A(state[1]), .B(state[0]), .Z(n2781)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_276.init = 16'h8888;
    LUT4 i5_4_lut (.A(state[3]), .B(n10_adj_198), .C(n22484), .D(state[1]), 
         .Z(n9453)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i5_4_lut.init = 16'h0040;
    LUT4 i4_4_lut_adj_277 (.A(\reset_count[14] ), .B(state[2]), .C(state[0]), 
         .D(n1156), .Z(n10_adj_198)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i4_4_lut_adj_277.init = 16'h0200;
    \ClockDividerP(factor=1250)  baud_gen (.GND_net(GND_net), .bclk(bclk), 
            .debug_c_c(debug_c_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=1250) 
//

module \ClockDividerP(factor=1250)  (GND_net, bclk, debug_c_c) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output bclk;
    input debug_c_c;
    
    wire bclk /* synthesis SET_AS_NETWORK=\motor_serial/sserial/sender/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27145;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n8542, n27144, n27143, n27142, n27141, n27140, n27139, 
        n27138, n27137, n27136, n27135, n27134, n27133, n27132, 
        n27131, n27067;
    wire [31:0]n102;
    
    wire n27066, n29844, n45, n52, n46, n16805, n50, n42, n27065, 
        n27064, n27063, n27062, n48, n38, n27061, n27060, n27059, 
        n44, n30, n29622, n27058, n27057, n27056, n27055, n27054, 
        n27053, n27052;
    
    CCU2D add_19626_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27145), 
          .S1(n8542));
    defparam add_19626_32.INIT0 = 16'h5555;
    defparam add_19626_32.INIT1 = 16'h0000;
    defparam add_19626_32.INJECT1_0 = "NO";
    defparam add_19626_32.INJECT1_1 = "NO";
    CCU2D add_19626_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27144), .COUT(n27145));
    defparam add_19626_30.INIT0 = 16'h5555;
    defparam add_19626_30.INIT1 = 16'h5555;
    defparam add_19626_30.INJECT1_0 = "NO";
    defparam add_19626_30.INJECT1_1 = "NO";
    CCU2D add_19626_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27143), .COUT(n27144));
    defparam add_19626_28.INIT0 = 16'h5555;
    defparam add_19626_28.INIT1 = 16'h5555;
    defparam add_19626_28.INJECT1_0 = "NO";
    defparam add_19626_28.INJECT1_1 = "NO";
    CCU2D add_19626_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27142), .COUT(n27143));
    defparam add_19626_26.INIT0 = 16'h5555;
    defparam add_19626_26.INIT1 = 16'h5555;
    defparam add_19626_26.INJECT1_0 = "NO";
    defparam add_19626_26.INJECT1_1 = "NO";
    CCU2D add_19626_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27141), .COUT(n27142));
    defparam add_19626_24.INIT0 = 16'h5555;
    defparam add_19626_24.INIT1 = 16'h5555;
    defparam add_19626_24.INJECT1_0 = "NO";
    defparam add_19626_24.INJECT1_1 = "NO";
    CCU2D add_19626_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27140), .COUT(n27141));
    defparam add_19626_22.INIT0 = 16'h5555;
    defparam add_19626_22.INIT1 = 16'h5555;
    defparam add_19626_22.INJECT1_0 = "NO";
    defparam add_19626_22.INJECT1_1 = "NO";
    CCU2D add_19626_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27139), .COUT(n27140));
    defparam add_19626_20.INIT0 = 16'h5555;
    defparam add_19626_20.INIT1 = 16'h5555;
    defparam add_19626_20.INJECT1_0 = "NO";
    defparam add_19626_20.INJECT1_1 = "NO";
    CCU2D add_19626_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27138), .COUT(n27139));
    defparam add_19626_18.INIT0 = 16'h5555;
    defparam add_19626_18.INIT1 = 16'h5555;
    defparam add_19626_18.INJECT1_0 = "NO";
    defparam add_19626_18.INJECT1_1 = "NO";
    CCU2D add_19626_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27137), .COUT(n27138));
    defparam add_19626_16.INIT0 = 16'h5555;
    defparam add_19626_16.INIT1 = 16'h5555;
    defparam add_19626_16.INJECT1_0 = "NO";
    defparam add_19626_16.INJECT1_1 = "NO";
    CCU2D add_19626_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27136), .COUT(n27137));
    defparam add_19626_14.INIT0 = 16'h5555;
    defparam add_19626_14.INIT1 = 16'h5555;
    defparam add_19626_14.INJECT1_0 = "NO";
    defparam add_19626_14.INJECT1_1 = "NO";
    CCU2D add_19626_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27135), .COUT(n27136));
    defparam add_19626_12.INIT0 = 16'h5555;
    defparam add_19626_12.INIT1 = 16'h5555;
    defparam add_19626_12.INJECT1_0 = "NO";
    defparam add_19626_12.INJECT1_1 = "NO";
    CCU2D add_19626_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27134), .COUT(n27135));
    defparam add_19626_10.INIT0 = 16'h5aaa;
    defparam add_19626_10.INIT1 = 16'h5555;
    defparam add_19626_10.INJECT1_0 = "NO";
    defparam add_19626_10.INJECT1_1 = "NO";
    CCU2D add_19626_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27133), 
          .COUT(n27134));
    defparam add_19626_8.INIT0 = 16'h5555;
    defparam add_19626_8.INIT1 = 16'h5555;
    defparam add_19626_8.INJECT1_0 = "NO";
    defparam add_19626_8.INJECT1_1 = "NO";
    CCU2D add_19626_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27132), 
          .COUT(n27133));
    defparam add_19626_6.INIT0 = 16'h5aaa;
    defparam add_19626_6.INIT1 = 16'h5aaa;
    defparam add_19626_6.INJECT1_0 = "NO";
    defparam add_19626_6.INJECT1_1 = "NO";
    CCU2D add_19626_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27131), 
          .COUT(n27132));
    defparam add_19626_4.INIT0 = 16'h5555;
    defparam add_19626_4.INIT1 = 16'h5aaa;
    defparam add_19626_4.INJECT1_0 = "NO";
    defparam add_19626_4.INJECT1_1 = "NO";
    CCU2D add_19626_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27131));
    defparam add_19626_2.INIT0 = 16'h1000;
    defparam add_19626_2.INIT1 = 16'h5555;
    defparam add_19626_2.INJECT1_0 = "NO";
    defparam add_19626_2.INJECT1_1 = "NO";
    FD1S3AX clk_o_14 (.D(n8542), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D count_2681_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27067), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_33.INIT1 = 16'h0000;
    defparam count_2681_add_4_33.INJECT1_0 = "NO";
    defparam count_2681_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2681_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27066), .COUT(n27067), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2681_add_4_31.INJECT1_0 = "NO";
    defparam count_2681_add_4_31.INJECT1_1 = "NO";
    LUT4 i22386_4_lut (.A(n29844), .B(n45), .C(n52), .D(n46), .Z(n16805)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i22386_4_lut.init = 16'h0002;
    LUT4 i22384_4_lut (.A(count[13]), .B(n50), .C(n42), .D(count[3]), 
         .Z(n29844)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i22384_4_lut.init = 16'h0001;
    LUT4 i17_4_lut (.A(count[26]), .B(count[12]), .C(count[9]), .D(count[17]), 
         .Z(n45)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i17_4_lut.init = 16'hfffe;
    CCU2D count_2681_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27065), .COUT(n27066), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2681_add_4_29.INJECT1_0 = "NO";
    defparam count_2681_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2681_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27064), .COUT(n27065), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2681_add_4_27.INJECT1_0 = "NO";
    defparam count_2681_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2681_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27063), .COUT(n27064), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2681_add_4_25.INJECT1_0 = "NO";
    defparam count_2681_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2681_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27062), .COUT(n27063), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2681_add_4_23.INJECT1_0 = "NO";
    defparam count_2681_add_4_23.INJECT1_1 = "NO";
    LUT4 i24_4_lut (.A(count[30]), .B(n48), .C(n38), .D(count[14]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(count[24]), .B(count[4]), .C(count[1]), .D(count[27]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i18_4_lut.init = 16'hfffe;
    CCU2D count_2681_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27061), .COUT(n27062), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2681_add_4_21.INJECT1_0 = "NO";
    defparam count_2681_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2681_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27060), .COUT(n27061), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2681_add_4_19.INJECT1_0 = "NO";
    defparam count_2681_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2681_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27059), .COUT(n27060), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2681_add_4_17.INJECT1_0 = "NO";
    defparam count_2681_add_4_17.INJECT1_1 = "NO";
    LUT4 i22_4_lut (.A(count[28]), .B(n44), .C(n30), .D(count[18]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(count[31]), .B(count[5]), .C(n29622), .D(count[6]), 
         .Z(n42)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i14_4_lut.init = 16'hbfff;
    CCU2D count_2681_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27058), .COUT(n27059), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2681_add_4_15.INJECT1_0 = "NO";
    defparam count_2681_add_4_15.INJECT1_1 = "NO";
    LUT4 i16_4_lut (.A(count[16]), .B(count[21]), .C(count[11]), .D(count[25]), 
         .Z(n44)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[2]), .B(count[8]), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(count[20]), .B(count[23]), .C(count[15]), .D(count[29]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i20_4_lut.init = 16'hfffe;
    CCU2D count_2681_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27057), .COUT(n27058), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2681_add_4_13.INJECT1_0 = "NO";
    defparam count_2681_add_4_13.INJECT1_1 = "NO";
    LUT4 i10_2_lut (.A(count[19]), .B(count[22]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i22063_3_lut (.A(count[10]), .B(count[0]), .C(count[7]), .Z(n29622)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i22063_3_lut.init = 16'h8080;
    CCU2D count_2681_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27056), .COUT(n27057), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2681_add_4_11.INJECT1_0 = "NO";
    defparam count_2681_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2681_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27055), .COUT(n27056), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2681_add_4_9.INJECT1_0 = "NO";
    defparam count_2681_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2681_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27054), .COUT(n27055), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2681_add_4_7.INJECT1_0 = "NO";
    defparam count_2681_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2681_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27053), .COUT(n27054), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2681_add_4_5.INJECT1_0 = "NO";
    defparam count_2681_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2681_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27052), .COUT(n27053), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2681_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2681_add_4_3.INJECT1_0 = "NO";
    defparam count_2681_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2681_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27052), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681_add_4_1.INIT0 = 16'hF000;
    defparam count_2681_add_4_1.INIT1 = 16'h0555;
    defparam count_2681_add_4_1.INJECT1_0 = "NO";
    defparam count_2681_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2681__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i0.GSR = "ENABLED";
    FD1S3IX count_2681__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i1.GSR = "ENABLED";
    FD1S3IX count_2681__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i2.GSR = "ENABLED";
    FD1S3IX count_2681__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i3.GSR = "ENABLED";
    FD1S3IX count_2681__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i4.GSR = "ENABLED";
    FD1S3IX count_2681__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i5.GSR = "ENABLED";
    FD1S3IX count_2681__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i6.GSR = "ENABLED";
    FD1S3IX count_2681__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i7.GSR = "ENABLED";
    FD1S3IX count_2681__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i8.GSR = "ENABLED";
    FD1S3IX count_2681__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i9.GSR = "ENABLED";
    FD1S3IX count_2681__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i10.GSR = "ENABLED";
    FD1S3IX count_2681__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i11.GSR = "ENABLED";
    FD1S3IX count_2681__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i12.GSR = "ENABLED";
    FD1S3IX count_2681__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i13.GSR = "ENABLED";
    FD1S3IX count_2681__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i14.GSR = "ENABLED";
    FD1S3IX count_2681__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i15.GSR = "ENABLED";
    FD1S3IX count_2681__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i16.GSR = "ENABLED";
    FD1S3IX count_2681__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i17.GSR = "ENABLED";
    FD1S3IX count_2681__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i18.GSR = "ENABLED";
    FD1S3IX count_2681__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i19.GSR = "ENABLED";
    FD1S3IX count_2681__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i20.GSR = "ENABLED";
    FD1S3IX count_2681__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i21.GSR = "ENABLED";
    FD1S3IX count_2681__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i22.GSR = "ENABLED";
    FD1S3IX count_2681__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i23.GSR = "ENABLED";
    FD1S3IX count_2681__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i24.GSR = "ENABLED";
    FD1S3IX count_2681__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i25.GSR = "ENABLED";
    FD1S3IX count_2681__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i26.GSR = "ENABLED";
    FD1S3IX count_2681__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i27.GSR = "ENABLED";
    FD1S3IX count_2681__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i28.GSR = "ENABLED";
    FD1S3IX count_2681__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i29.GSR = "ENABLED";
    FD1S3IX count_2681__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i30.GSR = "ENABLED";
    FD1S3IX count_2681__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n16805), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2681__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000) 
//

module \ClockDividerP(factor=12000)  (GND_net, n8507, n29786, n31512, 
            select_clk, \state[0] , n14037, n12, debug_c_c, n2967, 
            n107) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n8507;
    output n29786;
    input n31512;
    output select_clk;
    input \state[0] ;
    output n14037;
    output n12;
    input debug_c_c;
    input n2967;
    input n107;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27158;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n27157, n27156, n27155, n27154, n27153, n27152, n27151, 
        n27150, n27149, n27148, n27147, n27146, n27782, n15, n20, 
        n16, n27, n40, n36, n28, n18, n38, n32;
    wire [31:0]n134;
    
    wire n34, n24, n27051, n27050, n27049, n27048, n27047, n27046, 
        n27045, n27044, n27043, n27042, n27041, n27040, n27039, 
        n27038, n27037, n27036;
    
    CCU2D add_19625_28 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27158), 
          .S1(n8507));
    defparam add_19625_28.INIT0 = 16'h5555;
    defparam add_19625_28.INIT1 = 16'h0000;
    defparam add_19625_28.INJECT1_0 = "NO";
    defparam add_19625_28.INJECT1_1 = "NO";
    CCU2D add_19625_26 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27157), .COUT(n27158));
    defparam add_19625_26.INIT0 = 16'h5555;
    defparam add_19625_26.INIT1 = 16'h5555;
    defparam add_19625_26.INJECT1_0 = "NO";
    defparam add_19625_26.INJECT1_1 = "NO";
    CCU2D add_19625_24 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27156), .COUT(n27157));
    defparam add_19625_24.INIT0 = 16'h5555;
    defparam add_19625_24.INIT1 = 16'h5555;
    defparam add_19625_24.INJECT1_0 = "NO";
    defparam add_19625_24.INJECT1_1 = "NO";
    CCU2D add_19625_22 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27155), .COUT(n27156));
    defparam add_19625_22.INIT0 = 16'h5555;
    defparam add_19625_22.INIT1 = 16'h5555;
    defparam add_19625_22.INJECT1_0 = "NO";
    defparam add_19625_22.INJECT1_1 = "NO";
    CCU2D add_19625_20 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27154), .COUT(n27155));
    defparam add_19625_20.INIT0 = 16'h5555;
    defparam add_19625_20.INIT1 = 16'h5555;
    defparam add_19625_20.INJECT1_0 = "NO";
    defparam add_19625_20.INJECT1_1 = "NO";
    CCU2D add_19625_18 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27153), .COUT(n27154));
    defparam add_19625_18.INIT0 = 16'h5555;
    defparam add_19625_18.INIT1 = 16'h5555;
    defparam add_19625_18.INJECT1_0 = "NO";
    defparam add_19625_18.INJECT1_1 = "NO";
    CCU2D add_19625_16 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27152), .COUT(n27153));
    defparam add_19625_16.INIT0 = 16'h5555;
    defparam add_19625_16.INIT1 = 16'h5555;
    defparam add_19625_16.INJECT1_0 = "NO";
    defparam add_19625_16.INJECT1_1 = "NO";
    CCU2D add_19625_14 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27151), .COUT(n27152));
    defparam add_19625_14.INIT0 = 16'h5555;
    defparam add_19625_14.INIT1 = 16'h5555;
    defparam add_19625_14.INJECT1_0 = "NO";
    defparam add_19625_14.INJECT1_1 = "NO";
    CCU2D add_19625_12 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27150), .COUT(n27151));
    defparam add_19625_12.INIT0 = 16'h5555;
    defparam add_19625_12.INIT1 = 16'h5555;
    defparam add_19625_12.INJECT1_0 = "NO";
    defparam add_19625_12.INJECT1_1 = "NO";
    CCU2D add_19625_10 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27149), .COUT(n27150));
    defparam add_19625_10.INIT0 = 16'h5555;
    defparam add_19625_10.INIT1 = 16'h5555;
    defparam add_19625_10.INJECT1_0 = "NO";
    defparam add_19625_10.INJECT1_1 = "NO";
    CCU2D add_19625_8 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27148), .COUT(n27149));
    defparam add_19625_8.INIT0 = 16'h5555;
    defparam add_19625_8.INIT1 = 16'h5aaa;
    defparam add_19625_8.INJECT1_0 = "NO";
    defparam add_19625_8.INJECT1_1 = "NO";
    CCU2D add_19625_6 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27147), .COUT(n27148));
    defparam add_19625_6.INIT0 = 16'h5aaa;
    defparam add_19625_6.INIT1 = 16'h5aaa;
    defparam add_19625_6.INJECT1_0 = "NO";
    defparam add_19625_6.INJECT1_1 = "NO";
    CCU2D add_19625_4 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27146), 
          .COUT(n27147));
    defparam add_19625_4.INIT0 = 16'h5555;
    defparam add_19625_4.INIT1 = 16'h5aaa;
    defparam add_19625_4.INJECT1_0 = "NO";
    defparam add_19625_4.INJECT1_1 = "NO";
    CCU2D add_19625_2 (.A0(count[5]), .B0(count[4]), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27146));
    defparam add_19625_2.INIT0 = 16'h7000;
    defparam add_19625_2.INIT1 = 16'h5aaa;
    defparam add_19625_2.INJECT1_0 = "NO";
    defparam add_19625_2.INJECT1_1 = "NO";
    LUT4 i22326_4_lut (.A(n27782), .B(n15), .C(n20), .D(n16), .Z(n29786)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i22326_4_lut.init = 16'h4000;
    LUT4 i20_4_lut (.A(n27), .B(n40), .C(n36), .D(n28), .Z(n27782)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(count[11]), .B(count[10]), .Z(n15)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4_2_lut.init = 16'h8888;
    LUT4 i9_4_lut (.A(count[9]), .B(n18), .C(count[6]), .D(count[7]), 
         .Z(n20)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i9_4_lut.init = 16'h8000;
    LUT4 i5_2_lut (.A(count[1]), .B(count[4]), .Z(n16)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5_2_lut.init = 16'h8888;
    LUT4 i22357_2_lut_4_lut (.A(n31512), .B(select_clk), .C(n8507), .D(\state[0] ), 
         .Z(n14037)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(23[5] 33[8])
    defparam i22357_2_lut_4_lut.init = 16'h0010;
    LUT4 i5969_2_lut_4_lut (.A(n31512), .B(select_clk), .C(n8507), .D(\state[0] ), 
         .Z(n12)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(23[5] 33[8])
    defparam i5969_2_lut_4_lut.init = 16'hef10;
    LUT4 i6_2_lut (.A(count[28]), .B(count[12]), .Z(n27)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i19_4_lut (.A(count[5]), .B(n38), .C(n32), .D(count[20]), .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i15_4_lut (.A(count[8]), .B(count[25]), .C(count[15]), .D(count[26]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i15_4_lut.init = 16'hfffe;
    FD1S3IX count_2680__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2967), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i0.GSR = "ENABLED";
    LUT4 i7_2_lut (.A(count[17]), .B(count[24]), .Z(n28)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i7_4_lut (.A(count[13]), .B(count[2]), .C(count[3]), .D(count[0]), 
         .Z(n18)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i17_4_lut (.A(count[29]), .B(n34), .C(n24), .D(count[14]), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i11_3_lut (.A(count[22]), .B(count[21]), .C(count[31]), .Z(n32)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_3_lut.init = 16'hfefe;
    LUT4 i13_4_lut (.A(count[16]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[19]), .B(count[18]), .Z(n24)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i3_2_lut.init = 16'heeee;
    FD1S3AX clk_o_14 (.D(n107), .CK(debug_c_c), .Q(select_clk)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=25, LSE_RCOL=48, LSE_LLINE=21, LSE_RLINE=23 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D count_2680_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27051), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_33.INIT1 = 16'h0000;
    defparam count_2680_add_4_33.INJECT1_0 = "NO";
    defparam count_2680_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27050), .COUT(n27051), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_31.INJECT1_0 = "NO";
    defparam count_2680_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27049), .COUT(n27050), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_29.INJECT1_0 = "NO";
    defparam count_2680_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27048), .COUT(n27049), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_27.INJECT1_0 = "NO";
    defparam count_2680_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27047), .COUT(n27048), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_25.INJECT1_0 = "NO";
    defparam count_2680_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27046), .COUT(n27047), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_23.INJECT1_0 = "NO";
    defparam count_2680_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27045), .COUT(n27046), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_21.INJECT1_0 = "NO";
    defparam count_2680_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27044), .COUT(n27045), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_19.INJECT1_0 = "NO";
    defparam count_2680_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27043), .COUT(n27044), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_17.INJECT1_0 = "NO";
    defparam count_2680_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27042), .COUT(n27043), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_15.INJECT1_0 = "NO";
    defparam count_2680_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27041), .COUT(n27042), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_13.INJECT1_0 = "NO";
    defparam count_2680_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27040), .COUT(n27041), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_11.INJECT1_0 = "NO";
    defparam count_2680_add_4_11.INJECT1_1 = "NO";
    FD1S3IX count_2680__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2967), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i1.GSR = "ENABLED";
    CCU2D count_2680_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27039), .COUT(n27040), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_9.INJECT1_0 = "NO";
    defparam count_2680_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27038), .COUT(n27039), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_7.INJECT1_0 = "NO";
    defparam count_2680_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27037), .COUT(n27038), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_5.INJECT1_0 = "NO";
    defparam count_2680_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27036), .COUT(n27037), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2680_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2680_add_4_3.INJECT1_0 = "NO";
    defparam count_2680_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2680_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27036), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680_add_4_1.INIT0 = 16'hF000;
    defparam count_2680_add_4_1.INIT1 = 16'h0555;
    defparam count_2680_add_4_1.INJECT1_0 = "NO";
    defparam count_2680_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2680__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2967), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i2.GSR = "ENABLED";
    FD1S3IX count_2680__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2967), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i3.GSR = "ENABLED";
    FD1S3IX count_2680__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2967), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i4.GSR = "ENABLED";
    FD1S3IX count_2680__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2967), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i5.GSR = "ENABLED";
    FD1S3IX count_2680__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2967), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i6.GSR = "ENABLED";
    FD1S3IX count_2680__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2967), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i7.GSR = "ENABLED";
    FD1S3IX count_2680__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2967), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i8.GSR = "ENABLED";
    FD1S3IX count_2680__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2967), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i9.GSR = "ENABLED";
    FD1S3IX count_2680__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i10.GSR = "ENABLED";
    FD1S3IX count_2680__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i11.GSR = "ENABLED";
    FD1S3IX count_2680__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i12.GSR = "ENABLED";
    FD1S3IX count_2680__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i13.GSR = "ENABLED";
    FD1S3IX count_2680__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i14.GSR = "ENABLED";
    FD1S3IX count_2680__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i15.GSR = "ENABLED";
    FD1S3IX count_2680__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i16.GSR = "ENABLED";
    FD1S3IX count_2680__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i17.GSR = "ENABLED";
    FD1S3IX count_2680__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i18.GSR = "ENABLED";
    FD1S3IX count_2680__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i19.GSR = "ENABLED";
    FD1S3IX count_2680__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i20.GSR = "ENABLED";
    FD1S3IX count_2680__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i21.GSR = "ENABLED";
    FD1S3IX count_2680__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i22.GSR = "ENABLED";
    FD1S3IX count_2680__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i23.GSR = "ENABLED";
    FD1S3IX count_2680__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i24.GSR = "ENABLED";
    FD1S3IX count_2680__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i25.GSR = "ENABLED";
    FD1S3IX count_2680__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i26.GSR = "ENABLED";
    FD1S3IX count_2680__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i27.GSR = "ENABLED";
    FD1S3IX count_2680__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i28.GSR = "ENABLED";
    FD1S3IX count_2680__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i29.GSR = "ENABLED";
    FD1S3IX count_2680__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i30.GSR = "ENABLED";
    FD1S3IX count_2680__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2967), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2680__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ProtocolInterface(baud_div=12) 
//

module \ProtocolInterface(baud_div=12)  (register_addr, debug_c_c, databus, 
            \select[7] , n33390, \select[5] , \select[4] , \select[3] , 
            \select[2] , \select[1] , databus_out, n13834, \sendcount[1] , 
            n31556, n29301, n31533, n29200, debug_c_5, n31497, rw, 
            n31426, prev_select, n31428, n31596, n31470, n31466, 
            n31427, \register[1][19] , n59, n31501, \register[1][20] , 
            n57, \register[1][26] , n45, force_pause, \register[2] , 
            \register[1][0] , n97, n31504, prev_select_adj_5, n31512, 
            n13941, n1492, n29170, n29295, n29069, n29293, n31436, 
            n303, n56, n29294, n29066, n29056, n29053, n29065, 
            n29063, n29050, n224, n3922, n29052, n29054, n27752, 
            n29067, n29057, n29068, n29071, n29072, n27753, n29070, 
            n29058, n29059, n29064, n29060, n29258, n29062, n29055, 
            n29051, n29049, n29061, n29048, prev_select_adj_6, n2847, 
            n66, \register[0][2] , read_value, n33385, n2, n31465, 
            n2_adj_7, n2_adj_8, n2_adj_9, n2_adj_10, n31541, n31450, 
            n31478, n31471, n2_adj_11, n2_adj_12, n2_adj_13, n31474, 
            n2_adj_14, n2_adj_15, n2_adj_16, n2_adj_17, n2_adj_18, 
            n2_adj_19, n2_adj_20, n2_adj_21, n2_adj_22, n2_adj_23, 
            n3, n3_adj_24, n3_adj_25, n31590, n31477, n3_adj_26, 
            n3_adj_27, n3_adj_28, n3_adj_29, n3_adj_30, n2_adj_31, 
            n2_adj_32, n2_adj_33, n2_adj_34, n2_adj_35, n2_adj_36, 
            n31483, n14454, n9538, n35, n27465, n33384, n31446, 
            debug_c_7, \read_size[2] , n29235, n31445, n52, n31443, 
            n29237, n176, n31449, n31571, n16013, n31457, n31582, 
            n13908, n11236, n31435, n30306, n29221, n31526, n31420, 
            n30304, \control_reg[7] , n1, n31530, n31540, n13156, 
            n13, n18, n14, \reg_size[2] , n31588, n31591, n27442, 
            \control_reg[7]_adj_37 , n31601, n32, n4, n5834, prev_select_adj_38, 
            \reset_count[14] , n22484, n2870, n224_adj_91, n4095, 
            n31576, \read_value[7]_adj_71 , n2_adj_72, \read_value[5]_adj_73 , 
            n2_adj_74, n31473, \read_value[4]_adj_75 , n2_adj_76, \read_value[6]_adj_77 , 
            n2_adj_78, \read_value[3]_adj_79 , n2_adj_80, \read_value[2]_adj_81 , 
            n2_adj_82, \read_value[0]_adj_83 , n2_adj_84, n27445, n34, 
            n29257, n9331, n1486, \register[0][5] , expansion5_c, 
            \register[1][5] , debug_c_2, n1489, debug_c_3, n9379, 
            n29492, prev_select_adj_85, \steps_reg[7] , n11, debug_c_4, 
            n31502, n6006, \steps_reg[5] , n14_adj_86, \register[0][4] , 
            expansion4_out, \register[1][4] , timeout_pause, \steps_reg[6] , 
            n13_adj_87, \register[0][7] , n31537, clk_1Hz, signal_light_c, 
            \steps_reg[3] , n12, \control_reg[4] , \div_factor_reg[4] , 
            \steps_reg[4] , \control_reg[7]_adj_88 , n8636, n13948, 
            n12369, n9301, n14523, n4007, n31407, n27680, n27484, 
            n32_adj_89, n16765, n9, n9305, prev_select_adj_90, n16764, 
            n6003, n27428, n28827, n8654, \state[3] , \state[1] , 
            \state[0] , n1156, n73, \reset_count[7] , \reset_count[6] , 
            \reset_count[5] , n27250, uart_tx_c, GND_net, uart_rx_c) /* synthesis syn_module_defined=1 */ ;
    output [7:0]register_addr;
    input debug_c_c;
    input [31:0]databus;
    output \select[7] ;
    input n33390;
    output \select[5] ;
    output \select[4] ;
    output \select[3] ;
    output \select[2] ;
    output \select[1] ;
    output [31:0]databus_out;
    input n13834;
    output \sendcount[1] ;
    output n31556;
    output n29301;
    output n31533;
    output n29200;
    output debug_c_5;
    output n31497;
    output rw;
    output n31426;
    input prev_select;
    output n31428;
    output n31596;
    output n31470;
    output n31466;
    output n31427;
    input \register[1][19] ;
    output n59;
    input n31501;
    input \register[1][20] ;
    output n57;
    input \register[1][26] ;
    output n45;
    input force_pause;
    input [31:0]\register[2] ;
    input \register[1][0] ;
    output n97;
    output n31504;
    input prev_select_adj_5;
    input n31512;
    output n13941;
    output n1492;
    input n29170;
    output n29295;
    output n29069;
    output n29293;
    output n31436;
    output n303;
    output n56;
    output n29294;
    output n29066;
    output n29056;
    output n29053;
    output n29065;
    output n29063;
    output n29050;
    input [31:0]n224;
    output [31:0]n3922;
    output n29052;
    output n29054;
    output n27752;
    output n29067;
    output n29057;
    output n29068;
    output n29071;
    output n29072;
    output n27753;
    output n29070;
    output n29058;
    output n29059;
    output n29064;
    output n29060;
    output n29258;
    output n29062;
    output n29055;
    output n29051;
    output n29049;
    output n29061;
    output n29048;
    input prev_select_adj_6;
    output n2847;
    output n66;
    input \register[0][2] ;
    input [31:0]read_value;
    output n33385;
    output n2;
    output n31465;
    output n2_adj_7;
    output n2_adj_8;
    output n2_adj_9;
    output n2_adj_10;
    input n31541;
    output n31450;
    output n31478;
    output n31471;
    output n2_adj_11;
    output n2_adj_12;
    output n2_adj_13;
    output n31474;
    output n2_adj_14;
    output n2_adj_15;
    output n2_adj_16;
    output n2_adj_17;
    output n2_adj_18;
    output n2_adj_19;
    output n2_adj_20;
    output n2_adj_21;
    output n2_adj_22;
    output n2_adj_23;
    output n3;
    output n3_adj_24;
    output n3_adj_25;
    output n31590;
    output n31477;
    output n3_adj_26;
    output n3_adj_27;
    output n3_adj_28;
    output n3_adj_29;
    output n3_adj_30;
    output n2_adj_31;
    output n2_adj_32;
    output n2_adj_33;
    output n2_adj_34;
    output n2_adj_35;
    output n2_adj_36;
    output n31483;
    input n14454;
    output n9538;
    input n35;
    input n27465;
    input n33384;
    output n31446;
    output debug_c_7;
    input \read_size[2] ;
    output n29235;
    output n31445;
    output n52;
    output n31443;
    input n29237;
    output n176;
    output n31449;
    output n31571;
    output n16013;
    output n31457;
    input n31582;
    output n13908;
    output n11236;
    output n31435;
    output n30306;
    output n29221;
    output n31526;
    output n31420;
    output n30304;
    input \control_reg[7] ;
    output n1;
    output n31530;
    output n31540;
    input n13156;
    input n13;
    input n18;
    input n14;
    input \reg_size[2] ;
    input n31588;
    input n31591;
    input n27442;
    input \control_reg[7]_adj_37 ;
    output n31601;
    output n32;
    output n4;
    output n5834;
    input prev_select_adj_38;
    input \reset_count[14] ;
    input n22484;
    output n2870;
    input [31:0]n224_adj_91;
    output [31:0]n4095;
    output n31576;
    input \read_value[7]_adj_71 ;
    output n2_adj_72;
    input \read_value[5]_adj_73 ;
    output n2_adj_74;
    input n31473;
    input \read_value[4]_adj_75 ;
    output n2_adj_76;
    input \read_value[6]_adj_77 ;
    output n2_adj_78;
    input \read_value[3]_adj_79 ;
    output n2_adj_80;
    input \read_value[2]_adj_81 ;
    output n2_adj_82;
    input \read_value[0]_adj_83 ;
    output n2_adj_84;
    input n27445;
    output n34;
    output n29257;
    output n9331;
    output n1486;
    input \register[0][5] ;
    input expansion5_c;
    input \register[1][5] ;
    output debug_c_2;
    output n1489;
    output debug_c_3;
    output n9379;
    output n29492;
    input prev_select_adj_85;
    input \steps_reg[7] ;
    output n11;
    output debug_c_4;
    output n31502;
    output n6006;
    input \steps_reg[5] ;
    output n14_adj_86;
    input \register[0][4] ;
    input expansion4_out;
    input \register[1][4] ;
    input timeout_pause;
    input \steps_reg[6] ;
    output n13_adj_87;
    input \register[0][7] ;
    output n31537;
    input clk_1Hz;
    output signal_light_c;
    input \steps_reg[3] ;
    output n12;
    input \control_reg[4] ;
    input \div_factor_reg[4] ;
    input \steps_reg[4] ;
    input \control_reg[7]_adj_88 ;
    output n8636;
    output n13948;
    output n12369;
    output n9301;
    output n14523;
    output n4007;
    output n31407;
    output n27680;
    input n27484;
    output n32_adj_89;
    output n16765;
    input n9;
    output n9305;
    input prev_select_adj_90;
    output n16764;
    output n6003;
    output n27428;
    output n28827;
    output n8654;
    input \state[3] ;
    input \state[1] ;
    input \state[0] ;
    input n1156;
    output n73;
    input \reset_count[7] ;
    input \reset_count[6] ;
    input \reset_count[5] ;
    output n27250;
    output uart_tx_c;
    input GND_net;
    input uart_rx_c;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(455[15:21])
    wire n33384 /* synthesis nomerge= */ ;
    
    wire n2806;
    wire [7:0]\buffer[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]\buffer[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [31:0]n1474;
    wire [7:0]rx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(50[13:20])
    
    wire n29358, n5, n5_adj_39, n29022, n27598, n5_adj_40, n29023, 
        n27539;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    
    wire n31476;
    wire [4:0]n15;
    
    wire n15668, n5_adj_41, n29024, n27549, n31401, n31400, n31647, 
        n16686, n31644, n2808;
    wire [7:0]\buffer[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]\buffer[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]\buffer[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]esc_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(51[12:20])
    wire [7:0]n5825;
    wire [3:0]bufcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(46[12:20])
    
    wire n31611, n33381, n15680;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(52[12:19])
    
    wire n31469;
    wire [7:0]n2216;
    
    wire n15783, n30708, n5_adj_42, n29025, n27557;
    wire [7:0]\buffer[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n9472, n28593, n31448, n30824, n5_adj_43, n29028, n27525, 
        n31613, n31612, n31544, n31549, n10, n31554, n11_c, n11_adj_44, 
        n11_adj_45, n11_adj_46, n11_adj_47, n11_adj_48, n11_adj_49, 
        n11_adj_50, n31619, n31618, n31950, n31952, n2747, n16770, 
        n31622, n31621, n31625, n31624, n30303, n28917, n29390, 
        n31628, n31627, n31631, n31630, n15675, n1927, n31634, 
        n31633, n31646, n15671;
    wire [4:0]n17;
    
    wire n27682, n31637, n31636, n27434, n31640, n31639, n31609, 
        n31610, n31642, n31645, n9_adj_53, n31584, n31506, n31643, 
        n31424, n5_adj_54, n29026, n27505, n31451, n31542;
    wire [3:0]n1870;
    
    wire n31415, n31423, n31586, n31535, n4_c, n31623;
    wire [7:0]n9241;
    
    wire n4_adj_55, n31626, n29359, n4_adj_56, n31614, n4_adj_57, 
        n31632, n13490, n29205, n31487, n5_adj_58, n29029, n27473, 
        n31454, n14_c, n5_adj_59, n29032, n27533, n29019, n29256, 
        n29020, n29021, n5_adj_60, n29031, n27558, n31508, escape, 
        n10975, n30305, n5_adj_62, n29027, n27492, n4_adj_63, n31638, 
        n4_adj_64, n31635, n5_adj_65, n29033, n27556, n5_adj_69, 
        n29034, n27555, n2225, n29035, n29030, n5_adj_71, n27552, 
        n29036, n29037, n31545, n5_adj_77, n27551, n29361, n29038, 
        n31585, n31641, n30706, n30707, n5_adj_82, n27501, n7, 
        n30340, n29574, n38, n4_adj_85, n31629, n29039, n29040, 
        n29041, n29042, n29043, n29044, n29045, n5_adj_88, n27544, 
        n5_adj_89, n27534, n29046, n30823, n5_adj_95, n27427, n29015, 
        n5_adj_97, n27479, n29018, n29016, n5_adj_98, n27611, n29017, 
        n31553, n27626, n5_adj_102, n27497, n5_adj_103, n27514, 
        n29362, n5_adj_107, n27513, n31600, n57_adj_109, n31479, 
        n5_adj_110, n27477, n11_adj_111, n11_adj_112, n11_adj_113, 
        n11_adj_114, n5_adj_115, n27512, n31552, n11_adj_116, n11_adj_117, 
        n11_adj_118, n11_adj_119, n5_adj_120, n27511, send, n5_adj_121, 
        n27466, n31513, n1875, n31550, n31551, n9_adj_122, n5_adj_123, 
        n27506, n6, n5_adj_124, n27500, n31515, n7_adj_125, n31523, 
        n28667, n28659, n31539, n28617, n31524, n29277, n28, n29231, 
        n28615, n28619, n28621, n28663, n15679, n1_adj_126, n6_adj_127, 
        n28613, n28661, n15782, n31507, n28625, n28609, n28611, 
        n30341, n28587, n28623, n28607, n5_adj_130, n27602, n5_adj_131, 
        n27600, n15667, n16685, n27603, n31416, n13789, n31581, 
        n30342, n30734, n13_adj_151, busy, n11203, n19332;
    wire [7:0]register_addr_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    
    wire n12350, n79, n159, n8, n10_adj_157, n13042, n45_adj_163, 
        n112, n28900, n25, n19, n12_adj_172, n6_adj_173, n29163, 
        n28693, n16768, n13465, n12482, n29229, n1579, n1585, 
        n1586, n11217, n12348, n28605, n8_adj_182, n8_adj_185, n7_adj_186, 
        n29648, n29560, n29424, n30736;
    
    FD1P3AX reg_addr_i0_i0 (.D(\buffer[1] [0]), .SP(n2806), .CK(debug_c_c), 
            .Q(register_addr[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i0.GSR = "ENABLED";
    LUT4 select_2130_Select_18_i5_4_lut (.A(\buffer[2] [2]), .B(n1474[4]), 
         .C(rx_data[2]), .D(n29358), .Z(n5)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_18_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut (.A(databus[3]), .B(n5_adj_39), .C(n1474[13]), .D(n29022), 
         .Z(n27598)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut.init = 16'hffec;
    LUT4 select_2130_Select_19_i5_4_lut (.A(\buffer[2] [3]), .B(n1474[4]), 
         .C(rx_data[3]), .D(n29358), .Z(n5_adj_39)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_19_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_82 (.A(databus[4]), .B(n5_adj_40), .C(n1474[13]), 
         .D(n29023), .Z(n27539)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_82.init = 16'hffec;
    LUT4 select_2130_Select_20_i5_4_lut (.A(\buffer[2] [4]), .B(n1474[4]), 
         .C(rx_data[4]), .D(n29358), .Z(n5_adj_40)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_20_i5_4_lut.init = 16'h88c0;
    FD1P3AX sendcount__i0 (.D(n15[0]), .SP(n31476), .CK(debug_c_c), .Q(sendcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i0.GSR = "ENABLED";
    FD1S3IX select__i7 (.D(n15668), .CK(debug_c_c), .CD(n33390), .Q(\select[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i7.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_83 (.A(databus[5]), .B(n5_adj_41), .C(n1474[13]), 
         .D(n29024), .Z(n27549)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_83.init = 16'hffec;
    FD1S3IX select__i5 (.D(n31401), .CK(debug_c_c), .CD(n33390), .Q(\select[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i5.GSR = "ENABLED";
    FD1S3IX select__i4 (.D(n31400), .CK(debug_c_c), .CD(n33390), .Q(\select[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i4.GSR = "ENABLED";
    FD1S3IX select__i3 (.D(n31647), .CK(debug_c_c), .CD(n33390), .Q(\select[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i3.GSR = "ENABLED";
    FD1S3IX select__i2 (.D(n16686), .CK(debug_c_c), .CD(n33390), .Q(\select[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i2.GSR = "ENABLED";
    FD1S3IX select__i1 (.D(n31644), .CK(debug_c_c), .CD(n33390), .Q(\select[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i1.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i31 (.D(\buffer[5] [7]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i31.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i30 (.D(\buffer[5] [6]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i30.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i29 (.D(\buffer[5] [5]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i29.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i28 (.D(\buffer[5] [4]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i28.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i27 (.D(\buffer[5] [3]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i27.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i26 (.D(\buffer[5] [2]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i26.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i25 (.D(\buffer[5] [1]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i25.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i24 (.D(\buffer[5] [0]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i24.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i23 (.D(\buffer[4] [7]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i23.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i22 (.D(\buffer[4] [6]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i22.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i21 (.D(\buffer[4] [5]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i21.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i20 (.D(\buffer[4] [4]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i20.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i19 (.D(\buffer[4] [3]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i19.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i18 (.D(\buffer[4] [2]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i18.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i17 (.D(\buffer[4] [1]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i17.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i16 (.D(\buffer[4] [0]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i16.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i15 (.D(\buffer[3] [7]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i15.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i14 (.D(\buffer[3] [6]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i14.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i13 (.D(\buffer[3] [5]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i13.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i12 (.D(\buffer[3] [4]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i12.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i11 (.D(\buffer[3] [3]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i11.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i10 (.D(\buffer[3] [2]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i10.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i9 (.D(\buffer[3] [1]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i9.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i8 (.D(\buffer[3] [0]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i8.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i7 (.D(\buffer[2] [7]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i7.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i6 (.D(\buffer[2] [6]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i6.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i5 (.D(\buffer[2] [5]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i5.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i4 (.D(\buffer[2] [4]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i4.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i3 (.D(\buffer[2] [3]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i3.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i2 (.D(\buffer[2] [2]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i2.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i1 (.D(\buffer[2] [1]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i1.GSR = "ENABLED";
    LUT4 select_2130_Select_21_i5_4_lut (.A(\buffer[2] [5]), .B(n1474[4]), 
         .C(rx_data[5]), .D(n29358), .Z(n5_adj_41)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_21_i5_4_lut.init = 16'h88c0;
    FD1P3AX esc_data_i0_i4 (.D(n5825[4]), .SP(n13834), .CK(debug_c_c), 
            .Q(esc_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i4.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i2 (.D(n5825[2]), .SP(n13834), .CK(debug_c_c), 
            .Q(esc_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i2.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i1 (.D(n5825[1]), .SP(n13834), .CK(debug_c_c), 
            .Q(esc_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i1.GSR = "ENABLED";
    FD1S3IX bufcount__i3 (.D(n31611), .CK(debug_c_c), .CD(n33390), .Q(bufcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i3.GSR = "ENABLED";
    FD1S3IX bufcount__i2 (.D(n33381), .CK(debug_c_c), .CD(n33390), .Q(bufcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i2.GSR = "ENABLED";
    FD1S3IX bufcount__i1 (.D(n15680), .CK(debug_c_c), .CD(n33390), .Q(bufcount[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i1.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i4 (.D(n2216[4]), .SP(n31469), .CK(debug_c_c), 
            .Q(tx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n2216[3]), .SP(n31469), .CK(debug_c_c), 
            .Q(tx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i1 (.D(n2216[1]), .SP(n31469), .CK(debug_c_c), 
            .Q(tx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i0 (.D(n2216[0]), .SP(n31469), .CK(debug_c_c), 
            .Q(tx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    FD1S3IX bufcount__i0 (.D(n15783), .CK(debug_c_c), .CD(n33390), .Q(bufcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i0.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i0 (.D(n30708), .SP(n13834), .CK(debug_c_c), .Q(esc_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i0.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i0 (.D(\buffer[2] [0]), .SP(n2808), .CK(debug_c_c), 
            .Q(databus_out[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i0.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_84 (.A(databus[6]), .B(n5_adj_42), .C(n1474[13]), 
         .D(n29025), .Z(n27557)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_84.init = 16'hffec;
    FD1P3IX buffer_0___i1 (.D(n28593), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i1.GSR = "ENABLED";
    LUT4 select_2130_Select_22_i5_4_lut (.A(\buffer[2] [6]), .B(n1474[4]), 
         .C(rx_data[6]), .D(n29358), .Z(n5_adj_42)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_22_i5_4_lut.init = 16'h88c0;
    FD1P3IX sendcount__i4 (.D(n30824), .SP(n31476), .CD(n31448), .CK(debug_c_c), 
            .Q(sendcount[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i4.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_85 (.A(databus[7]), .B(n5_adj_43), .C(n1474[13]), 
         .D(n29028), .Z(n27525)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_85.init = 16'hffec;
    LUT4 i22192_then_3_lut (.A(\buffer[0] [5]), .B(\buffer[2] [5]), .C(\sendcount[1] ), 
         .Z(n31613)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22192_then_3_lut.init = 16'hcaca;
    LUT4 i22192_else_3_lut (.A(\buffer[3] [5]), .B(\buffer[1] [5]), .C(\sendcount[1] ), 
         .Z(n31612)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22192_else_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(register_addr[1]), .B(n31556), .C(register_addr[4]), 
         .D(n31544), .Z(n29301)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut.init = 16'h0002;
    LUT4 i2_2_lut_3_lut_4_lut (.A(register_addr[1]), .B(n31556), .C(n31533), 
         .D(register_addr[4]), .Z(n29200)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i5_3_lut_4_lut (.A(n31549), .B(n1474[12]), .C(n10), .D(n1474[9]), 
         .Z(debug_c_5)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5_3_lut_4_lut.init = 16'hfffe;
    LUT4 i24_3_lut_4_lut (.A(bufcount[0]), .B(n31554), .C(\buffer[0] [0]), 
         .D(rx_data[0]), .Z(n11_c)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_86 (.A(bufcount[0]), .B(n31554), .C(rx_data[1]), 
         .D(\buffer[0] [1]), .Z(n11_adj_44)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_86.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_87 (.A(bufcount[0]), .B(n31554), .C(rx_data[2]), 
         .D(\buffer[0] [2]), .Z(n11_adj_45)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_87.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_88 (.A(bufcount[0]), .B(n31554), .C(\buffer[0] [3]), 
         .D(rx_data[3]), .Z(n11_adj_46)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_88.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_89 (.A(bufcount[0]), .B(n31554), .C(\buffer[0] [4]), 
         .D(rx_data[4]), .Z(n11_adj_47)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_89.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_90 (.A(bufcount[0]), .B(n31554), .C(\buffer[0] [5]), 
         .D(rx_data[5]), .Z(n11_adj_48)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_90.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_91 (.A(bufcount[0]), .B(n31554), .C(\buffer[0] [6]), 
         .D(rx_data[6]), .Z(n11_adj_49)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_91.init = 16'hf1e0;
    LUT4 i20_2_lut_rep_282_3_lut_4_lut (.A(\select[4] ), .B(n31497), .C(rw), 
         .D(register_addr[5]), .Z(n31426)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i20_2_lut_rep_282_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_284_3_lut_4_lut (.A(\select[4] ), .B(n31497), .C(prev_select), 
         .D(register_addr[5]), .Z(n31428)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_284_3_lut_4_lut.init = 16'h0800;
    LUT4 i24_3_lut_4_lut_adj_92 (.A(bufcount[0]), .B(n31554), .C(rx_data[7]), 
         .D(\buffer[0] [7]), .Z(n11_adj_50)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_92.init = 16'hfe10;
    LUT4 i1_2_lut_rep_326_3_lut_4_lut (.A(register_addr[4]), .B(n31596), 
         .C(register_addr[5]), .D(n31556), .Z(n31470)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_2_lut_rep_326_3_lut_4_lut.init = 16'h0002;
    LUT4 i1_4_lut_then_4_lut (.A(sendcount[4]), .B(\sendcount[1] ), .C(sendcount[0]), 
         .D(sendcount[2]), .Z(n31619)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_rep_322_3_lut_4_lut (.A(register_addr[4]), .B(n31596), 
         .C(\select[4] ), .D(n31556), .Z(n31466)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_2_lut_rep_322_3_lut_4_lut.init = 16'h0020;
    LUT4 i1_4_lut_else_4_lut (.A(sendcount[4]), .B(\sendcount[1] ), .C(sendcount[0]), 
         .D(sendcount[2]), .Z(n31618)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h4001;
    LUT4 n31950_bdd_4_lut (.A(n31950), .B(n1474[4]), .C(n31952), .D(bufcount[2]), 
         .Z(n33381)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n31950_bdd_4_lut.init = 16'heef0;
    LUT4 i1_2_lut_3_lut (.A(register_addr[0]), .B(n31427), .C(\register[1][19] ), 
         .Z(n59)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i15753_3_lut_rep_325 (.A(n2747), .B(n31501), .C(n1474[18]), .Z(n31469)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i15753_3_lut_rep_325.init = 16'hc8c8;
    LUT4 i22347_2_lut_3_lut (.A(n2747), .B(n31501), .C(n1474[18]), .Z(n16770)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i22347_2_lut_3_lut.init = 16'h0808;
    LUT4 i22177_then_3_lut (.A(\buffer[0] [7]), .B(\buffer[2] [7]), .C(\sendcount[1] ), 
         .Z(n31622)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22177_then_3_lut.init = 16'hcaca;
    LUT4 i22177_else_3_lut (.A(\buffer[3] [7]), .B(\buffer[1] [7]), .C(\sendcount[1] ), 
         .Z(n31621)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22177_else_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_93 (.A(register_addr[0]), .B(n31427), .C(\register[1][20] ), 
         .Z(n57)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_adj_93.init = 16'h2020;
    LUT4 i22180_then_3_lut (.A(\buffer[0] [6]), .B(\buffer[2] [6]), .C(\sendcount[1] ), 
         .Z(n31625)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22180_then_3_lut.init = 16'hcaca;
    LUT4 i22180_else_3_lut (.A(\buffer[3] [6]), .B(\buffer[1] [6]), .C(\sendcount[1] ), 
         .Z(n31624)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22180_else_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_94 (.A(register_addr[0]), .B(n31427), .C(\register[1][26] ), 
         .Z(n45)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_adj_94.init = 16'h2020;
    LUT4 force_pause_bdd_4_lut (.A(force_pause), .B(register_addr[0]), .C(register_addr[1]), 
         .D(\register[2] [1]), .Z(n30303)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D))))) */ ;
    defparam force_pause_bdd_4_lut.init = 16'h3e0e;
    LUT4 i1_2_lut_3_lut_adj_95 (.A(register_addr[0]), .B(n31427), .C(\register[1][0] ), 
         .Z(n97)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_adj_95.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_96 (.A(\buffer[0] [1]), .B(n28917), .C(\buffer[0] [2]), 
         .Z(n29390)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i1_2_lut_3_lut_adj_96.init = 16'hefef;
    LUT4 i22195_then_3_lut (.A(\buffer[0] [4]), .B(\buffer[2] [4]), .C(\sendcount[1] ), 
         .Z(n31628)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22195_then_3_lut.init = 16'hcaca;
    LUT4 i22195_else_3_lut (.A(\buffer[3] [4]), .B(\buffer[1] [4]), .C(\sendcount[1] ), 
         .Z(n31627)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22195_else_3_lut.init = 16'hcaca;
    LUT4 i22198_then_3_lut (.A(\buffer[0] [3]), .B(\buffer[2] [3]), .C(\sendcount[1] ), 
         .Z(n31631)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22198_then_3_lut.init = 16'hcaca;
    LUT4 i22198_else_3_lut (.A(\buffer[3] [3]), .B(\buffer[1] [3]), .C(\sendcount[1] ), 
         .Z(n31630)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22198_else_3_lut.init = 16'hcaca;
    LUT4 \buffer_0[[0__bdd_4_lut_22979  (.A(\buffer[0] [0]), .B(n29390), 
         .C(n15675), .D(n1927), .Z(n31400)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;
    defparam \buffer_0[[0__bdd_4_lut_22979 .init = 16'h11f0;
    LUT4 i22201_then_3_lut (.A(\buffer[0] [2]), .B(\buffer[2] [2]), .C(\sendcount[1] ), 
         .Z(n31634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22201_then_3_lut.init = 16'hcaca;
    LUT4 i22201_else_3_lut (.A(\buffer[3] [2]), .B(\buffer[1] [2]), .C(\sendcount[1] ), 
         .Z(n31633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22201_else_3_lut.init = 16'hcaca;
    LUT4 n13751_bdd_4_lut_then_3_lut_4_lut (.A(\buffer[0] [2]), .B(\buffer[0] [0]), 
         .C(n28917), .D(\buffer[0] [1]), .Z(n31646)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam n13751_bdd_4_lut_then_3_lut_4_lut.init = 16'h0400;
    LUT4 \buffer_0[[0__bdd_4_lut  (.A(\buffer[0] [0]), .B(n29390), .C(n15671), 
         .D(n1927), .Z(n31401)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C))) */ ;
    defparam \buffer_0[[0__bdd_4_lut .init = 16'h22f0;
    FD1P3IX sendcount__i3 (.D(n17[3]), .SP(n31476), .CD(n31448), .CK(debug_c_c), 
            .Q(sendcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i3.GSR = "ENABLED";
    FD1P3IX sendcount__i2 (.D(n17[2]), .SP(n31476), .CD(n31448), .CK(debug_c_c), 
            .Q(sendcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i2.GSR = "ENABLED";
    FD1P3IX sendcount__i1 (.D(n17[1]), .SP(n31476), .CD(n31448), .CK(debug_c_c), 
            .Q(\sendcount[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i1.GSR = "ENABLED";
    LUT4 i22425_3_lut_4_lut (.A(\buffer[0] [1]), .B(n28917), .C(\buffer[0] [0]), 
         .D(\buffer[0] [2]), .Z(n27682)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i22425_3_lut_4_lut.init = 16'h2000;
    LUT4 i22204_then_3_lut (.A(\buffer[0] [1]), .B(\buffer[2] [1]), .C(\sendcount[1] ), 
         .Z(n31637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22204_then_3_lut.init = 16'hcaca;
    LUT4 i22204_else_3_lut (.A(\buffer[3] [1]), .B(\buffer[1] [1]), .C(\sendcount[1] ), 
         .Z(n31636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22204_else_3_lut.init = 16'hcaca;
    LUT4 i22465_3_lut_4_lut (.A(\buffer[0] [1]), .B(n28917), .C(\buffer[0] [0]), 
         .D(\buffer[0] [2]), .Z(n27434)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i22465_3_lut_4_lut.init = 16'h0002;
    LUT4 i22640_then_3_lut (.A(\buffer[0] [0]), .B(\buffer[2] [0]), .C(\sendcount[1] ), 
         .Z(n31640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22640_then_3_lut.init = 16'hcaca;
    LUT4 i22640_else_3_lut (.A(\buffer[3] [0]), .B(\buffer[1] [0]), .C(\sendcount[1] ), 
         .Z(n31639)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22640_else_3_lut.init = 16'hcaca;
    LUT4 i8898_else_4_lut (.A(bufcount[3]), .B(n1474[0]), .C(n1474[3]), 
         .D(n1474[4]), .Z(n31609)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i8898_else_4_lut.init = 16'h0002;
    LUT4 i8898_then_4_lut (.A(bufcount[3]), .B(n1474[0]), .C(n1474[3]), 
         .D(n1474[4]), .Z(n31610)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i8898_then_4_lut.init = 16'haaa2;
    LUT4 n13674_bdd_4_lut_else_3_lut (.A(\select[1] ), .B(n1474[8]), .C(n1474[0]), 
         .Z(n31642)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam n13674_bdd_4_lut_else_3_lut.init = 16'h0202;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(\select[4] ), .B(n31504), .C(prev_select_adj_5), 
         .D(n31512), .Z(n13941)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 n13751_bdd_4_lut_else_3_lut (.A(\select[3] ), .B(n1474[8]), .C(n1474[0]), 
         .Z(n31645)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam n13751_bdd_4_lut_else_3_lut.init = 16'h0202;
    LUT4 i15751_3_lut_rep_332 (.A(n1474[13]), .B(n31501), .C(n1492), .Z(n31476)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i15751_3_lut_rep_332.init = 16'hc8c8;
    LUT4 i14817_4_lut (.A(sendcount[3]), .B(n9_adj_53), .C(sendcount[2]), 
         .D(n31584), .Z(n17[3])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(271[10:37])
    defparam i14817_4_lut.init = 16'h4888;
    LUT4 i22350_2_lut_rep_304_3_lut (.A(n1474[13]), .B(n31501), .C(n1492), 
         .Z(n31448)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i22350_2_lut_rep_304_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_3_lut_4_lut (.A(register_addr[2]), .B(n31506), .C(\register[2] [31]), 
         .D(n29170), .Z(n29295)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_97 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [28]), .D(n29170), .Z(n29069)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_97.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_98 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [29]), .D(n29170), .Z(n29293)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_98.init = 16'h1000;
    LUT4 select_2130_Select_23_i5_4_lut (.A(\buffer[2] [7]), .B(n1474[4]), 
         .C(rx_data[7]), .D(n29358), .Z(n5_adj_43)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_23_i5_4_lut.init = 16'h88c0;
    LUT4 n13674_bdd_4_lut_then_3_lut_4_lut (.A(\buffer[0] [2]), .B(\buffer[0] [0]), 
         .C(n28917), .D(\buffer[0] [1]), .Z(n31643)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam n13674_bdd_4_lut_then_3_lut_4_lut.init = 16'h0004;
    LUT4 register_addr_1__bdd_3_lut_22612_rep_292_4_lut (.A(register_addr[2]), 
         .B(n31506), .C(register_addr[0]), .D(register_addr[1]), .Z(n31436)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam register_addr_1__bdd_3_lut_22612_rep_292_4_lut.init = 16'h0110;
    LUT4 i21972_2_lut_rep_280_3_lut_4_lut (.A(register_addr[2]), .B(n31506), 
         .C(rw), .D(register_addr[1]), .Z(n31424)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i21972_2_lut_rep_280_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_99 (.A(register_addr[2]), .B(n31506), 
         .C(register_addr[0]), .D(register_addr[1]), .Z(n303)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_99.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_4_lut_adj_100 (.A(register_addr[2]), .B(n31506), 
         .C(register_addr[0]), .D(register_addr[1]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_100.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_101 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [30]), .D(n29170), .Z(n29294)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_101.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_102 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [4]), .D(n29170), .Z(n29066)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_102.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_103 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [5]), .D(n29170), .Z(n29056)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_103.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_104 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [6]), .D(n29170), .Z(n29053)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_104.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_105 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [7]), .D(n29170), .Z(n29065)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_105.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_106 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [8]), .D(n29170), .Z(n29063)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_106.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_107 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [9]), .D(n29170), .Z(n29050)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_107.init = 16'h1000;
    LUT4 i2_4_lut_adj_108 (.A(databus[8]), .B(n5_adj_54), .C(n1474[13]), 
         .D(n29026), .Z(n27505)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_108.init = 16'hffec;
    LUT4 i3352_2_lut_3_lut_4_lut_4_lut (.A(bufcount[1]), .B(n31451), .C(n31542), 
         .D(bufcount[0]), .Z(n1870[1])) /* synthesis lut_function=(A (B (C+!(D)))+!A !((C+!(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i3352_2_lut_3_lut_4_lut_4_lut.init = 16'h8488;
    LUT4 mux_1554_i13_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[12]), 
         .D(n224[12]), .Z(n3922[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_109 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [10]), .D(n29170), .Z(n29052)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_109.init = 16'h1000;
    LUT4 mux_429_Mux_7_i7_4_lut_4_lut (.A(n31586), .B(n31535), .C(n4_c), 
         .D(n31623), .Z(n9241[7])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_7_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_6_i7_4_lut_4_lut (.A(n31586), .B(n31535), .C(n4_adj_55), 
         .D(n31626), .Z(n9241[6])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_6_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 select_2130_Select_24_i5_4_lut (.A(\buffer[3] [0]), .B(n1474[4]), 
         .C(rx_data[0]), .D(n29359), .Z(n5_adj_54)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_24_i5_4_lut.init = 16'h88c0;
    LUT4 mux_429_Mux_5_i7_4_lut_4_lut (.A(n31586), .B(n31535), .C(n4_adj_56), 
         .D(n31614), .Z(n9241[5])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_5_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_3_i7_4_lut_4_lut (.A(n31586), .B(n31535), .C(n4_adj_57), 
         .D(n31632), .Z(n9241[3])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_3_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i1_2_lut_3_lut_4_lut_adj_110 (.A(n31554), .B(bufcount[3]), .C(\buffer[0] [7]), 
         .D(n13490), .Z(n29205)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_110.init = 16'h0e00;
    LUT4 i22114_2_lut_rep_343_4_lut (.A(register_addr[5]), .B(n31596), .C(register_addr[4]), 
         .D(n31556), .Z(n31487)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22114_2_lut_rep_343_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_111 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [11]), .D(n29170), .Z(n29054)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_111.init = 16'h1000;
    LUT4 i22342_3_lut_4_lut (.A(n31556), .B(register_addr[1]), .C(register_addr[4]), 
         .D(n31533), .Z(n27752)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i22342_3_lut_4_lut.init = 16'h0010;
    LUT4 i2_4_lut_adj_112 (.A(databus[9]), .B(n5_adj_58), .C(n1474[13]), 
         .D(n29029), .Z(n27473)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_112.init = 16'hffec;
    LUT4 i1_2_lut_3_lut_4_lut_adj_113 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [12]), .D(n29170), .Z(n29067)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_113.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_114 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [13]), .D(n29170), .Z(n29057)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_114.init = 16'h1000;
    LUT4 select_2130_Select_25_i5_4_lut (.A(\buffer[3] [1]), .B(n1474[4]), 
         .C(rx_data[1]), .D(n29359), .Z(n5_adj_58)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_25_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_115 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [14]), .D(n29170), .Z(n29068)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_115.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_116 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [15]), .D(n29170), .Z(n29071)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_116.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_adj_117 (.A(n1474[3]), .B(n31454), .C(n1474[13]), 
         .Z(n14_c)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_117.init = 16'hf8f8;
    LUT4 i1_2_lut_3_lut_4_lut_adj_118 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [16]), .D(n29170), .Z(n29072)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_118.init = 16'h1000;
    LUT4 i22339_3_lut_4_lut (.A(n31556), .B(register_addr[1]), .C(register_addr[4]), 
         .D(n31544), .Z(n27753)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i22339_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_4_lut_adj_119 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [17]), .D(n29170), .Z(n29070)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_119.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_120 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [18]), .D(n29170), .Z(n29058)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_120.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_121 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [19]), .D(n29170), .Z(n29059)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_121.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_122 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [20]), .D(n29170), .Z(n29064)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_122.init = 16'h1000;
    LUT4 i2_4_lut_adj_123 (.A(databus[10]), .B(n5_adj_59), .C(n1474[13]), 
         .D(n29032), .Z(n27533)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_123.init = 16'hffec;
    LUT4 i1_2_lut_3_lut_4_lut_adj_124 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [21]), .D(n29170), .Z(n29060)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_124.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_adj_125 (.A(n1474[3]), .B(n31454), .C(\buffer[2] [0]), 
         .Z(n29019)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_125.init = 16'h8080;
    LUT4 select_2130_Select_26_i5_4_lut (.A(\buffer[3] [2]), .B(n1474[4]), 
         .C(rx_data[2]), .D(n29359), .Z(n5_adj_59)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_26_i5_4_lut.init = 16'h88c0;
    LUT4 i1_3_lut_4_lut (.A(n31556), .B(register_addr[1]), .C(n29256), 
         .D(n31596), .Z(n29258)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_4_lut_adj_126 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [22]), .D(n29170), .Z(n29062)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_126.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_adj_127 (.A(n1474[3]), .B(n31454), .C(\buffer[2] [1]), 
         .Z(n29020)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_127.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_128 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [23]), .D(n29170), .Z(n29055)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_128.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_129 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [24]), .D(n29170), .Z(n29051)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_129.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_adj_130 (.A(n1474[3]), .B(n31454), .C(\buffer[2] [2]), 
         .Z(n29021)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_130.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_131 (.A(n1474[3]), .B(n31454), .C(\buffer[2] [3]), 
         .Z(n29022)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_131.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_132 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [25]), .D(n29170), .Z(n29049)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_132.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_133 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [26]), .D(n29170), .Z(n29061)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_133.init = 16'h1000;
    FD1P3AX rw_498 (.D(n1474[10]), .SP(n2806), .CK(debug_c_c), .Q(rw));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_134 (.A(n1474[3]), .B(n31454), .C(\buffer[2] [4]), 
         .Z(n29023)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_134.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_135 (.A(register_addr[2]), .B(n31506), 
         .C(\register[2] [27]), .D(n29170), .Z(n29048)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_135.init = 16'h1000;
    LUT4 i2_4_lut_adj_136 (.A(databus[11]), .B(n5_adj_60), .C(n1474[13]), 
         .D(n29031), .Z(n27558)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_136.init = 16'hffec;
    LUT4 i1_2_lut_3_lut_adj_137 (.A(n1474[3]), .B(n31454), .C(\buffer[2] [5]), 
         .Z(n29024)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_137.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_138 (.A(n31508), .B(prev_select_adj_6), 
         .C(\select[4] ), .D(n31512), .Z(n2847)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_138.init = 16'h0010;
    LUT4 i1_2_lut (.A(\select[5] ), .B(rw), .Z(n66)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(454[7:9])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_139 (.A(n1474[3]), .B(n31454), .C(\buffer[2] [6]), 
         .Z(n29025)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_139.init = 16'h8080;
    FD1S3AX escape_501 (.D(n10975), .CK(debug_c_c), .Q(escape));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam escape_501.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_140 (.A(n1474[3]), .B(n31454), .C(\buffer[2] [7]), 
         .Z(n29028)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_140.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_141 (.A(n1474[3]), .B(n31454), .C(\buffer[3] [0]), 
         .Z(n29026)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_141.init = 16'h8080;
    LUT4 select_2130_Select_27_i5_4_lut (.A(\buffer[3] [3]), .B(n1474[4]), 
         .C(rx_data[3]), .D(n29359), .Z(n5_adj_60)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_27_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_142 (.A(n1474[3]), .B(n31454), .C(\buffer[3] [1]), 
         .Z(n29029)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_142.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_143 (.A(n1474[3]), .B(n31454), .C(\buffer[3] [2]), 
         .Z(n29032)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_143.init = 16'h8080;
    LUT4 \register_0[[2__bdd_4_lut  (.A(\register[0][2] ), .B(register_addr[0]), 
         .C(register_addr[1]), .D(\register[2] [2]), .Z(n30305)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D))))) */ ;
    defparam \register_0[[2__bdd_4_lut .init = 16'h3e0e;
    LUT4 i2_4_lut_adj_144 (.A(databus[12]), .B(n5_adj_62), .C(n1474[13]), 
         .D(n29027), .Z(n27492)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_144.init = 16'hffec;
    LUT4 mux_429_Mux_1_i7_4_lut_4_lut (.A(n31586), .B(n31535), .C(n4_adj_63), 
         .D(n31638), .Z(n9241[1])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_1_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 select_2130_Select_28_i5_4_lut (.A(\buffer[3] [4]), .B(n1474[4]), 
         .C(rx_data[4]), .D(n29359), .Z(n5_adj_62)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_28_i5_4_lut.init = 16'h88c0;
    LUT4 mux_429_Mux_2_i7_4_lut_4_lut (.A(n31586), .B(n31535), .C(n4_adj_64), 
         .D(n31635), .Z(n9241[2])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_2_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i1_2_lut_3_lut_adj_145 (.A(n1474[3]), .B(n31454), .C(\buffer[3] [3]), 
         .Z(n29031)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_145.init = 16'h8080;
    LUT4 Select_4244_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[23]), .D(n33385), .Z(n2)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4244_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_146 (.A(n1474[3]), .B(n31454), .C(\buffer[3] [4]), 
         .Z(n29027)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_146.init = 16'h8080;
    LUT4 i2_4_lut_adj_147 (.A(databus[13]), .B(n5_adj_65), .C(n1474[13]), 
         .D(n29033), .Z(n27556)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_147.init = 16'hffec;
    LUT4 select_2130_Select_29_i5_4_lut (.A(\buffer[3] [5]), .B(n1474[4]), 
         .C(rx_data[5]), .D(n29359), .Z(n5_adj_65)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_29_i5_4_lut.init = 16'h88c0;
    LUT4 i14703_2_lut_rep_321_3_lut_4_lut (.A(register_addr[5]), .B(n31596), 
         .C(\select[3] ), .D(register_addr[4]), .Z(n31465)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i14703_2_lut_rep_321_3_lut_4_lut.init = 16'he0f0;
    LUT4 Select_4247_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[22]), .D(n33385), .Z(n2_adj_7)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4247_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4250_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[21]), .D(n33385), .Z(n2_adj_8)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4250_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4253_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[20]), .D(n33385), .Z(n2_adj_9)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4253_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_148 (.A(n1474[3]), .B(n31454), .C(\buffer[3] [5]), 
         .Z(n29033)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_148.init = 16'h8080;
    LUT4 i2_4_lut_adj_149 (.A(databus[14]), .B(n5_adj_69), .C(n1474[13]), 
         .D(n29034), .Z(n27555)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_149.init = 16'hffec;
    LUT4 Select_4238_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[25]), .D(rw), .Z(n2_adj_10)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4238_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i22_1_lut_rep_306_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31596), 
         .C(n31541), .D(register_addr[4]), .Z(n31450)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i22_1_lut_rep_306_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_adj_150 (.A(n1474[3]), .B(n31454), .C(\buffer[3] [6]), 
         .Z(n29034)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_150.init = 16'h8080;
    LUT4 i1_2_lut_adj_151 (.A(n1474[16]), .B(n1474[19]), .Z(n2225)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_151.init = 16'heeee;
    LUT4 select_2130_Select_30_i5_4_lut (.A(\buffer[3] [6]), .B(n1474[4]), 
         .C(rx_data[6]), .D(n29359), .Z(n5_adj_69)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_30_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_152 (.A(n1474[3]), .B(n31454), .C(\buffer[3] [7]), 
         .Z(n29035)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_152.init = 16'h8080;
    LUT4 i1_2_lut_rep_334_3_lut_4_lut (.A(register_addr[5]), .B(n31596), 
         .C(n31541), .D(register_addr[4]), .Z(n31478)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_334_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_153 (.A(n1474[3]), .B(n31454), .C(\buffer[4] [0]), 
         .Z(n29030)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_153.init = 16'h8080;
    LUT4 i2_4_lut_adj_154 (.A(databus[15]), .B(n5_adj_71), .C(n1474[13]), 
         .D(n29035), .Z(n27552)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_154.init = 16'hffec;
    LUT4 i15037_2_lut_rep_327_3_lut_4_lut (.A(register_addr[5]), .B(n31596), 
         .C(\select[3] ), .D(register_addr[4]), .Z(n31471)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i15037_2_lut_rep_327_3_lut_4_lut.init = 16'h1000;
    LUT4 select_2130_Select_31_i5_4_lut (.A(\buffer[3] [7]), .B(n1474[4]), 
         .C(rx_data[7]), .D(n29359), .Z(n5_adj_71)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_31_i5_4_lut.init = 16'h88c0;
    LUT4 Select_4241_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[24]), .D(n33385), .Z(n2_adj_11)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4241_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4256_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[19]), .D(n33385), .Z(n2_adj_12)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4256_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_155 (.A(n1474[3]), .B(n31454), .C(\buffer[4] [1]), 
         .Z(n29036)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_155.init = 16'h8080;
    LUT4 Select_4259_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[18]), .D(rw), .Z(n2_adj_13)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4259_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_156 (.A(n1474[3]), .B(n31454), .C(\buffer[4] [2]), 
         .Z(n29037)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_156.init = 16'h8080;
    LUT4 i1_2_lut_rep_330_3_lut_4_lut (.A(register_addr[5]), .B(n31596), 
         .C(\select[4] ), .D(n31545), .Z(n31474)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_330_3_lut_4_lut.init = 16'h0010;
    LUT4 Select_4262_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[17]), .D(rw), .Z(n2_adj_14)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4262_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4265_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[16]), .D(rw), .Z(n2_adj_15)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4265_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_adj_157 (.A(databus[16]), .B(n5_adj_77), .C(n1474[13]), 
         .D(n29030), .Z(n27551)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_157.init = 16'hffec;
    LUT4 select_2130_Select_32_i5_4_lut (.A(\buffer[4] [0]), .B(n1474[4]), 
         .C(rx_data[0]), .D(n29361), .Z(n5_adj_77)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_32_i5_4_lut.init = 16'h88c0;
    LUT4 Select_4268_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[15]), .D(rw), .Z(n2_adj_16)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4268_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4271_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[14]), .D(rw), .Z(n2_adj_17)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4271_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_158 (.A(n1474[3]), .B(n31454), .C(\buffer[4] [3]), 
         .Z(n29038)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_158.init = 16'h8080;
    LUT4 Select_4274_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[13]), .D(rw), .Z(n2_adj_18)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4274_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 n30706_bdd_3_lut_4_lut (.A(sendcount[2]), .B(n31585), .C(n31641), 
         .D(n30706), .Z(n30707)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam n30706_bdd_3_lut_4_lut.init = 16'hf960;
    LUT4 Select_4277_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[12]), .D(rw), .Z(n2_adj_19)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4277_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_adj_159 (.A(databus[17]), .B(n5_adj_82), .C(n1474[13]), 
         .D(n29036), .Z(n27501)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_159.init = 16'hffec;
    LUT4 select_2130_Select_33_i5_4_lut (.A(\buffer[4] [1]), .B(n1474[4]), 
         .C(rx_data[1]), .D(n29361), .Z(n5_adj_82)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_33_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut (.A(n1474[15]), .B(n7), .C(n30340), .D(n29574), .Z(n38)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut.init = 16'haaa8;
    LUT4 Select_4280_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[11]), .D(rw), .Z(n2_adj_20)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4280_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4283_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[10]), .D(rw), .Z(n2_adj_21)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4283_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 mux_429_Mux_4_i7_4_lut_4_lut (.A(n31586), .B(n31535), .C(n4_adj_85), 
         .D(n31629), .Z(n9241[4])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_4_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i1_2_lut_3_lut_adj_160 (.A(n1474[3]), .B(n31454), .C(\buffer[4] [4]), 
         .Z(n29039)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_160.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_161 (.A(n1474[3]), .B(n31454), .C(\buffer[4] [5]), 
         .Z(n29040)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_161.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_162 (.A(n1474[3]), .B(n31454), .C(\buffer[4] [6]), 
         .Z(n29041)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_162.init = 16'h8080;
    LUT4 Select_4286_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[9]), .D(rw), .Z(n2_adj_22)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4286_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4289_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[8]), .D(rw), .Z(n2_adj_23)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4289_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_163 (.A(n1474[3]), .B(n31454), .C(\buffer[4] [7]), 
         .Z(n29042)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_163.init = 16'h8080;
    LUT4 Select_4290_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[7]), .D(rw), .Z(n3)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4290_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_164 (.A(n1474[3]), .B(n31454), .C(\buffer[5] [0]), 
         .Z(n29043)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_164.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_165 (.A(n1474[3]), .B(n31454), .C(\buffer[5] [1]), 
         .Z(n29044)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_165.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_166 (.A(n1474[3]), .B(n31454), .C(\buffer[5] [2]), 
         .Z(n29045)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_166.init = 16'h8080;
    LUT4 i2_4_lut_adj_167 (.A(databus[18]), .B(n5_adj_88), .C(n1474[13]), 
         .D(n29037), .Z(n27544)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_167.init = 16'hffec;
    LUT4 select_2130_Select_34_i5_4_lut (.A(\buffer[4] [2]), .B(n1474[4]), 
         .C(rx_data[2]), .D(n29361), .Z(n5_adj_88)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_34_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_168 (.A(databus[19]), .B(n5_adj_89), .C(n1474[13]), 
         .D(n29038), .Z(n27534)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_168.init = 16'hffec;
    LUT4 Select_4291_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[6]), .D(rw), .Z(n3_adj_24)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4291_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4292_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[5]), .D(rw), .Z(n3_adj_25)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4292_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_169 (.A(n1474[3]), .B(n31454), .C(\buffer[5] [3]), 
         .Z(n29046)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_169.init = 16'h8080;
    LUT4 sendcount_1__bdd_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(sendcount[3]), 
         .D(sendcount[2]), .Z(n30823)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;
    defparam sendcount_1__bdd_4_lut.init = 16'h6aaa;
    LUT4 select_2130_Select_35_i5_4_lut (.A(\buffer[4] [3]), .B(n1474[4]), 
         .C(rx_data[3]), .D(n29361), .Z(n5_adj_89)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_35_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_333_3_lut_4_lut (.A(register_addr[3]), .B(n31596), 
         .C(register_addr[2]), .D(n31590), .Z(n31477)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_333_3_lut_4_lut.init = 16'hfffe;
    LUT4 Select_4293_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[4]), .D(rw), .Z(n3_adj_26)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4293_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4294_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[3]), .D(rw), .Z(n3_adj_27)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4294_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4295_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[2]), .D(rw), .Z(n3_adj_28)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4295_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_adj_170 (.A(databus[20]), .B(n5_adj_95), .C(n1474[13]), 
         .D(n29039), .Z(n27427)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_170.init = 16'hffec;
    LUT4 Select_4296_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[1]), .D(rw), .Z(n3_adj_29)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4296_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 select_2130_Select_36_i5_4_lut (.A(\buffer[4] [4]), .B(n1474[4]), 
         .C(rx_data[4]), .D(n29361), .Z(n5_adj_95)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_36_i5_4_lut.init = 16'h88c0;
    LUT4 sendcount_4__bdd_3_lut (.A(sendcount[4]), .B(n30823), .C(\sendcount[1] ), 
         .Z(n30824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam sendcount_4__bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_171 (.A(n1474[3]), .B(n31454), .C(\buffer[5] [4]), 
         .Z(n29015)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_171.init = 16'h8080;
    LUT4 i2_4_lut_adj_172 (.A(databus[21]), .B(n5_adj_97), .C(n1474[13]), 
         .D(n29040), .Z(n27479)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_172.init = 16'hffec;
    LUT4 select_2130_Select_37_i5_4_lut (.A(\buffer[4] [5]), .B(n1474[4]), 
         .C(rx_data[5]), .D(n29361), .Z(n5_adj_97)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_37_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_173 (.A(n1474[3]), .B(n31454), .C(\buffer[5] [5]), 
         .Z(n29018)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_173.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_174 (.A(n1474[3]), .B(n31454), .C(\buffer[5] [6]), 
         .Z(n29016)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_174.init = 16'h8080;
    LUT4 i2_4_lut_adj_175 (.A(databus[22]), .B(n5_adj_98), .C(n1474[13]), 
         .D(n29041), .Z(n27611)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_175.init = 16'hffec;
    LUT4 Select_4297_i3_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[0]), .D(rw), .Z(n3_adj_30)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4297_i3_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 select_2130_Select_38_i5_4_lut (.A(\buffer[4] [6]), .B(n1474[4]), 
         .C(rx_data[6]), .D(n29361), .Z(n5_adj_98)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_38_i5_4_lut.init = 16'h88c0;
    LUT4 Select_4220_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[31]), .D(rw), .Z(n2_adj_31)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4220_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_176 (.A(n1474[3]), .B(n31454), .C(\buffer[5] [7]), 
         .Z(n29017)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_176.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_adj_177 (.A(n1474[4]), .B(n31553), .C(bufcount[0]), 
         .D(n31451), .Z(n27626)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_adj_177.init = 16'hd222;
    LUT4 Select_4223_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[30]), .D(rw), .Z(n2_adj_32)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4223_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_adj_178 (.A(databus[23]), .B(n5_adj_102), .C(n1474[13]), 
         .D(n29042), .Z(n27497)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_178.init = 16'hffec;
    LUT4 select_2130_Select_39_i5_4_lut (.A(\buffer[4] [7]), .B(n1474[4]), 
         .C(rx_data[7]), .D(n29361), .Z(n5_adj_102)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_39_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_179 (.A(databus[24]), .B(n5_adj_103), .C(n1474[13]), 
         .D(n29043), .Z(n27514)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_179.init = 16'hffec;
    LUT4 select_2130_Select_40_i5_4_lut (.A(\buffer[5] [0]), .B(n1474[4]), 
         .C(rx_data[0]), .D(n29362), .Z(n5_adj_103)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_40_i5_4_lut.init = 16'h88c0;
    LUT4 Select_4226_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[29]), .D(rw), .Z(n2_adj_33)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4226_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4229_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[28]), .D(rw), .Z(n2_adj_34)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4229_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4232_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[27]), .D(rw), .Z(n2_adj_35)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4232_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_adj_180 (.A(databus[25]), .B(n5_adj_107), .C(n1474[13]), 
         .D(n29044), .Z(n27513)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_180.init = 16'hffec;
    LUT4 Select_4235_i2_2_lut_3_lut_4_lut (.A(\select[4] ), .B(n31508), 
         .C(read_value[26]), .D(rw), .Z(n2_adj_36)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4235_i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i17816_3_lut_4_lut (.A(n31501), .B(n31600), .C(n57_adj_109), 
         .D(escape), .Z(n10975)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i17816_3_lut_4_lut.init = 16'h7780;
    LUT4 select_2130_Select_41_i5_4_lut (.A(\buffer[5] [1]), .B(n1474[4]), 
         .C(rx_data[1]), .D(n29362), .Z(n5_adj_107)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_41_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_335_3_lut_4_lut (.A(n31596), .B(register_addr[5]), 
         .C(prev_select_adj_6), .D(n31545), .Z(n31479)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_2_lut_rep_335_3_lut_4_lut.init = 16'hfffb;
    LUT4 mux_1554_i12_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[11]), 
         .D(n224[11]), .Z(n3922[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_339_3_lut_4_lut (.A(n31596), .B(register_addr[5]), 
         .C(\select[4] ), .D(n31545), .Z(n31483)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_rep_339_3_lut_4_lut.init = 16'h0040;
    LUT4 mux_1554_i19_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[18]), 
         .D(n224[18]), .Z(n3922[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1554_i18_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[17]), 
         .D(n224[17]), .Z(n3922[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_4_lut_adj_181 (.A(databus[26]), .B(n5_adj_110), .C(n1474[13]), 
         .D(n29045), .Z(n27477)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_181.init = 16'hffec;
    LUT4 i1_2_lut_rep_360_3_lut_4_lut (.A(register_addr[4]), .B(n31556), 
         .C(n31596), .D(register_addr[5]), .Z(n31504)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_360_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_364_3_lut_4_lut (.A(register_addr[4]), .B(n31556), 
         .C(register_addr[5]), .D(n31596), .Z(n31508)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_364_3_lut_4_lut.init = 16'hffef;
    LUT4 select_2130_Select_42_i5_4_lut (.A(\buffer[5] [2]), .B(n1474[4]), 
         .C(rx_data[2]), .D(n29362), .Z(n5_adj_110)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_42_i5_4_lut.init = 16'h88c0;
    LUT4 i24_3_lut_4_lut_adj_182 (.A(bufcount[0]), .B(n31554), .C(\buffer[1] [0]), 
         .D(rx_data[0]), .Z(n11_adj_111)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_182.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_183 (.A(bufcount[0]), .B(n31554), .C(rx_data[1]), 
         .D(\buffer[1] [1]), .Z(n11_adj_112)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_183.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_184 (.A(bufcount[0]), .B(n31554), .C(rx_data[2]), 
         .D(\buffer[1] [2]), .Z(n11_adj_113)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_184.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_185 (.A(bufcount[0]), .B(n31554), .C(\buffer[1] [3]), 
         .D(rx_data[3]), .Z(n11_adj_114)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_185.init = 16'hf2d0;
    LUT4 i2_4_lut_adj_186 (.A(databus[27]), .B(n5_adj_115), .C(n1474[13]), 
         .D(n29046), .Z(n27512)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_186.init = 16'hffec;
    LUT4 i2_3_lut_4_lut_adj_187 (.A(register_addr[1]), .B(n31477), .C(register_addr[0]), 
         .D(n14454), .Z(n9538)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut_adj_187.init = 16'h2000;
    LUT4 n31454_bdd_4_lut_23120 (.A(n31454), .B(n31552), .C(n1474[0]), 
         .D(n1474[3]), .Z(n31950)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam n31454_bdd_4_lut_23120.init = 16'hee0f;
    LUT4 i24_3_lut_4_lut_adj_188 (.A(bufcount[0]), .B(n31554), .C(\buffer[1] [4]), 
         .D(rx_data[4]), .Z(n11_adj_116)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_188.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_189 (.A(bufcount[0]), .B(n31554), .C(\buffer[1] [5]), 
         .D(rx_data[5]), .Z(n11_adj_117)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_189.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_190 (.A(bufcount[0]), .B(n31554), .C(rx_data[6]), 
         .D(\buffer[1] [6]), .Z(n11_adj_118)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_190.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_191 (.A(bufcount[0]), .B(n31554), .C(\buffer[1] [7]), 
         .D(rx_data[7]), .Z(n11_adj_119)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_191.init = 16'hf2d0;
    LUT4 select_2130_Select_43_i5_4_lut (.A(\buffer[5] [3]), .B(n1474[4]), 
         .C(rx_data[3]), .D(n29362), .Z(n5_adj_115)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_43_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_279 (.A(register_addr[4]), .B(n35), .Z(n31423)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_279.init = 16'h8888;
    LUT4 mux_1554_i17_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[16]), 
         .D(n224[16]), .Z(n3922[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_4_lut_adj_192 (.A(databus[28]), .B(n5_adj_120), .C(n1474[13]), 
         .D(n29015), .Z(n27511)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_192.init = 16'hffec;
    FD1P3IX send_491 (.D(n33384), .SP(n2225), .CD(n27465), .CK(debug_c_c), 
            .Q(send));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam send_491.GSR = "ENABLED";
    LUT4 select_2130_Select_44_i5_4_lut (.A(\buffer[5] [4]), .B(n1474[4]), 
         .C(rx_data[4]), .D(n29362), .Z(n5_adj_120)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_44_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_193 (.A(databus[29]), .B(n5_adj_121), .C(n1474[13]), 
         .D(n29018), .Z(n27466)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_193.init = 16'hffec;
    LUT4 i4_2_lut_rep_405 (.A(n1492), .B(n1474[15]), .Z(n31549)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_2_lut_rep_405.init = 16'heeee;
    LUT4 select_2130_Select_45_i5_4_lut (.A(\buffer[5] [5]), .B(n1474[4]), 
         .C(rx_data[5]), .D(n29362), .Z(n5_adj_121)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_45_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_369_3_lut (.A(n1492), .B(n1474[15]), .C(n1474[12]), 
         .Z(n31513)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_369_3_lut.init = 16'hfefe;
    LUT4 i508_2_lut (.A(n1474[3]), .B(n1474[4]), .Z(n1875)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i508_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_rep_406 (.A(n1474[19]), .B(n1474[3]), .C(n1474[11]), 
         .Z(n31550)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_3_lut_rep_406.init = 16'hfefe;
    LUT4 i3_2_lut_4_lut (.A(n1474[19]), .B(n1474[3]), .C(n1474[11]), .D(n31551), 
         .Z(n9_adj_122)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_2_lut_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_194 (.A(databus[30]), .B(n5_adj_123), .C(n1474[13]), 
         .D(n29016), .Z(n27506)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_194.init = 16'hffec;
    LUT4 select_2130_Select_46_i5_4_lut (.A(\buffer[5] [6]), .B(n1474[4]), 
         .C(rx_data[6]), .D(n29362), .Z(n5_adj_123)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_46_i5_4_lut.init = 16'h88c0;
    LUT4 i2_3_lut_rep_407 (.A(n1474[7]), .B(n1474[13]), .C(n1474[5]), 
         .Z(n31551)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_407.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut (.A(n1474[7]), .B(n1474[13]), .C(n1474[5]), .D(n1474[6]), 
         .Z(n6)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    LUT4 mux_1554_i11_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[10]), 
         .D(n224[10]), .Z(n3922[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_4_lut_adj_195 (.A(databus[31]), .B(n5_adj_124), .C(n1474[13]), 
         .D(n29017), .Z(n27500)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_195.init = 16'hffec;
    LUT4 select_2130_Select_47_i5_4_lut (.A(\buffer[5] [7]), .B(n1474[4]), 
         .C(rx_data[7]), .D(n29362), .Z(n5_adj_124)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_47_i5_4_lut.init = 16'h88c0;
    LUT4 n31454_bdd_4_lut (.A(bufcount[1]), .B(n1474[4]), .C(bufcount[0]), 
         .D(bufcount[3]), .Z(n31952)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam n31454_bdd_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_302_3_lut_4_lut (.A(n31556), .B(n31515), .C(\select[4] ), 
         .D(register_addr[5]), .Z(n31446)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_302_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_408 (.A(debug_c_7), .B(escape), .Z(n31552)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut_rep_408.init = 16'hdddd;
    LUT4 i2_3_lut_rep_307_4_lut (.A(debug_c_7), .B(escape), .C(n31454), 
         .D(n1474[4]), .Z(n31451)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i2_3_lut_rep_307_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_3_lut_4_lut_adj_196 (.A(n31556), .B(n31515), .C(\read_size[2] ), 
         .D(register_addr[5]), .Z(n29235)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_196.init = 16'h0040;
    LUT4 i1_2_lut_rep_301_3_lut_4_lut (.A(n31556), .B(n31515), .C(register_addr[5]), 
         .D(\select[4] ), .Z(n31445)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_301_3_lut_4_lut.init = 16'h4000;
    LUT4 i15597_3_lut_rep_409 (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .Z(n31553)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i15597_3_lut_rep_409.init = 16'hecec;
    LUT4 i2_2_lut_rep_398_4_lut (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1474[4]), .Z(n31542)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+!(D))) */ ;
    defparam i2_2_lut_rep_398_4_lut.init = 16'hecff;
    LUT4 i1_2_lut_4_lut_adj_197 (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1474[4]), .Z(n7_adj_125)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i1_2_lut_4_lut_adj_197.init = 16'hec00;
    LUT4 equal_202_i4_2_lut_rep_410 (.A(bufcount[1]), .B(bufcount[2]), .Z(n31554)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam equal_202_i4_2_lut_rep_410.init = 16'heeee;
    LUT4 mux_1554_i16_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[15]), 
         .D(n224[15]), .Z(n3922[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1554_i15_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[14]), 
         .D(n224[14]), .Z(n3922[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 i2938_2_lut_rep_379_3_lut (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[3]), 
         .Z(n31523)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i2938_2_lut_rep_379_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_198 (.A(n31545), .B(n31533), .C(n33385), 
         .D(\select[4] ), .Z(n52)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_198.init = 16'h1000;
    LUT4 i1_4_lut_adj_199 (.A(n1474[4]), .B(\buffer[0] [1]), .C(n11_adj_44), 
         .D(n14_c), .Z(n28667)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_199.init = 16'heca0;
    LUT4 i1_4_lut_adj_200 (.A(n1474[4]), .B(\buffer[0] [2]), .C(n11_adj_45), 
         .D(n14_c), .Z(n28659)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_200.init = 16'heca0;
    LUT4 i1_2_lut_rep_299_3_lut_4_lut (.A(n31545), .B(n31533), .C(prev_select_adj_5), 
         .D(\select[4] ), .Z(n31443)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_299_3_lut_4_lut.init = 16'h0100;
    LUT4 mux_1554_i14_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[13]), 
         .D(n224[13]), .Z(n3922[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i15592_1_lut_3_lut_4_lut (.A(n31590), .B(n31539), .C(n29237), 
         .D(register_addr[2]), .Z(n176)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i15592_1_lut_3_lut_4_lut.init = 16'h0111;
    LUT4 i1_2_lut_3_lut_4_lut_adj_201 (.A(rw), .B(n31449), .C(register_addr[0]), 
         .D(n31571), .Z(n16013)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_201.init = 16'h1000;
    LUT4 i15591_3_lut_rep_313_4_lut (.A(n31590), .B(n31539), .C(n29237), 
         .D(register_addr[2]), .Z(n31457)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i15591_3_lut_rep_313_4_lut.init = 16'hfeee;
    LUT4 i22018_2_lut (.A(esc_data[5]), .B(esc_data[6]), .Z(n29574)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22018_2_lut.init = 16'heeee;
    LUT4 i22361_2_lut_3_lut_4_lut (.A(rw), .B(n31449), .C(register_addr[0]), 
         .D(n31582), .Z(n13908)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i22361_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i21902_2_lut_rep_412 (.A(register_addr[2]), .B(register_addr[3]), 
         .Z(n31556)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21902_2_lut_rep_412.init = 16'heeee;
    LUT4 i4461_2_lut_3_lut_4_lut (.A(rw), .B(n31449), .C(register_addr[0]), 
         .D(n31582), .Z(n11236)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i4461_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_291_3_lut_4_lut (.A(n31590), .B(n31539), .C(register_addr[1]), 
         .D(register_addr[2]), .Z(n31435)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_291_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_4_lut_adj_202 (.A(n1474[4]), .B(\buffer[0] [3]), .C(n11_adj_46), 
         .D(n14_c), .Z(n28617)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_202.init = 16'heca0;
    LUT4 n30305_bdd_2_lut_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(n30305), .D(n31524), .Z(n30306)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam n30305_bdd_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 mux_1554_i10_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[9]), 
         .D(n224[9]), .Z(n3922[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 esc_data_1__bdd_4_lut (.A(esc_data[1]), .B(esc_data[3]), .C(esc_data[2]), 
         .D(esc_data[4]), .Z(n30340)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C (D)))+!A (B+(C+(D)))) */ ;
    defparam esc_data_1__bdd_4_lut.init = 16'hd7fe;
    LUT4 i1_2_lut_adj_203 (.A(rx_data[4]), .B(rx_data[1]), .Z(n29277)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_203.init = 16'h8888;
    LUT4 mux_1554_i1_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[0]), 
         .D(n224[0]), .Z(n3922[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1554_i32_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[31]), 
         .D(n224[31]), .Z(n3922[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i32_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_3_lut_4_lut_adj_204 (.A(register_addr[2]), .B(register_addr[3]), 
         .C(n28), .D(n31524), .Z(n29221)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_3_lut_4_lut_adj_204.init = 16'h0010;
    LUT4 mux_1554_i31_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[30]), 
         .D(n224[30]), .Z(n3922[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i31_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_305_3_lut_4_lut (.A(n31590), .B(n31539), .C(register_addr[1]), 
         .D(register_addr[2]), .Z(n31449)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_305_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21963_2_lut_rep_382_3_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[1]), .Z(n31526)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i21963_2_lut_rep_382_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_276_3_lut_4_lut (.A(register_addr[4]), .B(n31541), 
         .C(n29231), .D(n31596), .Z(n31420)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_276_3_lut_4_lut.init = 16'h0010;
    LUT4 n30303_bdd_2_lut_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(n30303), .D(n31524), .Z(n30304)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam n30303_bdd_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_adj_205 (.A(register_addr[0]), .B(\control_reg[7] ), .Z(n1)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_205.init = 16'h4444;
    LUT4 i1_4_lut_adj_206 (.A(n1474[4]), .B(\buffer[0] [4]), .C(n11_adj_47), 
         .D(n14_c), .Z(n28615)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_206.init = 16'heca0;
    LUT4 i2_3_lut_rep_386_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(n31596), .D(n29170), .Z(n31530)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_3_lut_rep_386_4_lut.init = 16'h0100;
    LUT4 i1_4_lut_adj_207 (.A(n1474[4]), .B(\buffer[0] [5]), .C(n11_adj_48), 
         .D(n14_c), .Z(n28619)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_207.init = 16'heca0;
    LUT4 i1_4_lut_adj_208 (.A(n1474[4]), .B(\buffer[0] [6]), .C(n11_adj_49), 
         .D(n14_c), .Z(n28621)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_208.init = 16'heca0;
    LUT4 i1_4_lut_adj_209 (.A(n1474[4]), .B(\buffer[0] [7]), .C(n11_adj_50), 
         .D(n14_c), .Z(n28663)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_209.init = 16'heca0;
    LUT4 i1_2_lut_rep_396_3_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[4]), .Z(n31540)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_396_3_lut.init = 16'h1010;
    PFUMX i8908 (.BLUT(n15679), .ALUT(n1870[1]), .C0(n1875), .Z(n15680));
    LUT4 i1_4_lut_adj_210 (.A(sendcount[4]), .B(n1_adj_126), .C(n6_adj_127), 
         .D(n13156), .Z(n9_adj_53)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i1_4_lut_adj_210.init = 16'hfeff;
    LUT4 equal_64_i1_4_lut (.A(sendcount[0]), .B(n13), .C(n18), .D(n14), 
         .Z(n1_adj_126)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam equal_64_i1_4_lut.init = 16'h5556;
    LUT4 i1_4_lut_adj_211 (.A(n1474[4]), .B(\buffer[1] [0]), .C(n11_adj_111), 
         .D(n14_c), .Z(n28613)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_211.init = 16'heca0;
    LUT4 i14917_2_lut (.A(bufcount[1]), .B(n1474[0]), .Z(n15679)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14917_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_212 (.A(\reg_size[2] ), .B(sendcount[3]), .C(sendcount[2]), 
         .D(n31588), .Z(n6_adj_127)) /* synthesis lut_function=(A (B (C+!(D))+!B ((D)+!C))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i2_4_lut_adj_212.init = 16'he7de;
    LUT4 i1_2_lut_3_lut_4_lut_adj_213 (.A(register_addr[2]), .B(register_addr[3]), 
         .C(n31596), .D(register_addr[4]), .Z(n31497)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_213.init = 16'h0100;
    LUT4 i1_4_lut_adj_214 (.A(n1474[4]), .B(\buffer[1] [1]), .C(n11_adj_112), 
         .D(n14_c), .Z(n28661)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_214.init = 16'heca0;
    PFUMX i9011 (.BLUT(n15782), .ALUT(n27626), .C0(n1875), .Z(n15783));
    LUT4 i1_2_lut_rep_363_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[4]), .D(n31591), .Z(n31507)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_363_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_215 (.A(n1474[4]), .B(\buffer[1] [2]), .C(n11_adj_113), 
         .D(n14_c), .Z(n28625)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_215.init = 16'heca0;
    LUT4 i1_2_lut_rep_401_3_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[4]), .Z(n31545)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_401_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_216 (.A(n1474[4]), .B(\buffer[1] [3]), .C(n11_adj_114), 
         .D(n14_c), .Z(n28609)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_216.init = 16'heca0;
    LUT4 i1_4_lut_adj_217 (.A(n1474[4]), .B(\buffer[1] [4]), .C(n11_adj_116), 
         .D(n14_c), .Z(n28611)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_217.init = 16'heca0;
    LUT4 n29162_bdd_4_lut (.A(sendcount[3]), .B(sendcount[2]), .C(sendcount[0]), 
         .D(\sendcount[1] ), .Z(n30341)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam n29162_bdd_4_lut.init = 16'h4001;
    LUT4 mux_1554_i30_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[29]), 
         .D(n224[29]), .Z(n3922[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i30_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_218 (.A(n1474[4]), .B(\buffer[1] [5]), .C(n11_adj_117), 
         .D(n14_c), .Z(n28587)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_218.init = 16'heca0;
    LUT4 i1_4_lut_adj_219 (.A(n1474[4]), .B(\buffer[1] [6]), .C(n11_adj_118), 
         .D(n14_c), .Z(n28623)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_219.init = 16'heca0;
    LUT4 mux_1554_i29_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[28]), 
         .D(n224[28]), .Z(n3922[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i29_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_220 (.A(n1474[4]), .B(\buffer[1] [7]), .C(n11_adj_119), 
         .D(n14_c), .Z(n28607)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_220.init = 16'heca0;
    LUT4 i2_4_lut_adj_221 (.A(databus[0]), .B(n5_adj_130), .C(n1474[13]), 
         .D(n29019), .Z(n27602)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_221.init = 16'hffec;
    LUT4 select_2130_Select_16_i5_4_lut (.A(\buffer[2] [0]), .B(n1474[4]), 
         .C(rx_data[0]), .D(n29358), .Z(n5_adj_130)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_16_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_222 (.A(databus[1]), .B(n5_adj_131), .C(n1474[13]), 
         .D(n29020), .Z(n27600)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_222.init = 16'hffec;
    LUT4 mux_1554_i9_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[8]), 
         .D(n224[8]), .Z(n3922[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1554_i28_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[27]), 
         .D(n224[27]), .Z(n3922[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i28_3_lut_4_lut.init = 16'hf780;
    LUT4 select_2130_Select_17_i5_4_lut (.A(\buffer[2] [1]), .B(n1474[4]), 
         .C(rx_data[1]), .D(n29358), .Z(n5_adj_131)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2130_Select_17_i5_4_lut.init = 16'h88c0;
    LUT4 i14922_2_lut_3_lut (.A(n1474[0]), .B(n1474[8]), .C(\select[7] ), 
         .Z(n15667)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i14922_2_lut_3_lut.init = 16'h1010;
    LUT4 i2_3_lut (.A(n27442), .B(\control_reg[7]_adj_37 ), .C(n31601), 
         .Z(n32)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut.init = 16'h0808;
    LUT4 mux_1554_i8_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[7]), 
         .D(n224[7]), .Z(n3922[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 i14920_2_lut_3_lut (.A(n1474[0]), .B(n1474[8]), .C(\select[5] ), 
         .Z(n15671)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i14920_2_lut_3_lut.init = 16'h1010;
    LUT4 i958_2_lut (.A(n1474[5]), .B(n31501), .Z(n2808)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i958_2_lut.init = 16'h8888;
    LUT4 i15120_2_lut_3_lut (.A(n1474[0]), .B(n1474[8]), .C(\select[2] ), 
         .Z(n16685)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i15120_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_223 (.A(n1474[0]), .B(n1474[8]), .C(\select[4] ), 
         .Z(n15675)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_223.init = 16'h1010;
    LUT4 i1_2_lut_adj_224 (.A(sendcount[0]), .B(sendcount[3]), .Z(n4)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_224.init = 16'h4444;
    LUT4 i2_4_lut_adj_225 (.A(databus[2]), .B(n5), .C(n1474[13]), .D(n29021), 
         .Z(n27603)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_225.init = 16'hffec;
    LUT4 mux_1896_i5_3_lut (.A(n9241[4]), .B(sendcount[0]), .C(n5834), 
         .Z(n5825[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1896_i5_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_4_i4_3_lut (.A(\buffer[4] [4]), .B(\buffer[5] [4]), 
         .C(sendcount[0]), .Z(n4_adj_85)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_4_i4_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_rep_427 (.A(\select[5] ), .B(prev_select_adj_38), .Z(n31571)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_427.init = 16'h2222;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(\select[5] ), .B(prev_select_adj_38), 
         .C(\reset_count[14] ), .D(n22484), .Z(n2870)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 mux_1554_i7_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[6]), 
         .D(n224[6]), .Z(n3922[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1554_i6_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[5]), 
         .D(n224[5]), .Z(n3922[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1599_i8_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[7]), 
         .D(n224_adj_91[7]), .Z(n4095[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1599_i7_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[6]), 
         .D(n224_adj_91[6]), .Z(n4095[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 i14930_2_lut (.A(bufcount[0]), .B(n1474[0]), .Z(n15782)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14930_2_lut.init = 16'h2222;
    LUT4 mux_1554_i5_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[4]), 
         .D(n224[4]), .Z(n3922[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1554_i4_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[3]), 
         .D(n224[3]), .Z(n3922[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_432 (.A(rw), .B(register_addr[5]), .Z(n31576)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_432.init = 16'h4444;
    LUT4 i1_2_lut_rep_271_3_lut_4_lut_4_lut (.A(n33385), .B(register_addr[5]), 
         .C(prev_select), .D(n31466), .Z(n31415)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_271_3_lut_4_lut_4_lut.init = 16'h0400;
    LUT4 Select_4290_i2_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31466), 
         .C(\read_value[7]_adj_71 ), .D(n33385), .Z(n2_adj_72)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4290_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_1896_i3_3_lut (.A(n9241[2]), .B(sendcount[0]), .C(n5834), 
         .Z(n5825[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1896_i3_3_lut.init = 16'hcaca;
    LUT4 Select_4292_i2_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31466), 
         .C(\read_value[5]_adj_73 ), .D(rw), .Z(n2_adj_74)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4292_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1S3JX state_FSM_i1 (.D(n13789), .CK(debug_c_c), .PD(n31473), .Q(n1474[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i1.GSR = "ENABLED";
    LUT4 mux_429_Mux_2_i4_3_lut (.A(\buffer[4] [2]), .B(\buffer[5] [2]), 
         .C(sendcount[0]), .Z(n4_adj_64)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_2_i4_3_lut.init = 16'hacac;
    LUT4 i956_3_lut (.A(n1474[5]), .B(n31501), .C(n1474[10]), .Z(n2806)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i956_3_lut.init = 16'hc8c8;
    LUT4 mux_1896_i2_3_lut (.A(n9241[1]), .B(sendcount[0]), .C(n5834), 
         .Z(n5825[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1896_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_437 (.A(n1492), .B(sendcount[4]), .Z(n31581)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_437.init = 16'h2222;
    LUT4 n1_bdd_2_lut_22586_3_lut (.A(n1492), .B(sendcount[4]), .C(n30341), 
         .Z(n30342)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam n1_bdd_2_lut_22586_3_lut.init = 16'h2020;
    LUT4 Select_4293_i2_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31466), 
         .C(\read_value[4]_adj_75 ), .D(rw), .Z(n2_adj_76)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4293_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_429_Mux_1_i4_3_lut (.A(\buffer[4] [1]), .B(\buffer[5] [1]), 
         .C(sendcount[0]), .Z(n4_adj_63)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_1_i4_3_lut.init = 16'hacac;
    PFUMX i9914 (.BLUT(n16685), .ALUT(n27434), .C0(n1927), .Z(n16686));
    PFUMX i8896 (.BLUT(n15667), .ALUT(n27682), .C0(n1927), .Z(n15668));
    LUT4 mux_1599_i20_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[19]), 
         .D(n224_adj_91[19]), .Z(n4095[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_522_i5_3_lut (.A(n2747), .B(esc_data[4]), .C(n1474[18]), 
         .Z(n2216[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_522_i5_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_226 (.A(n1474[15]), .B(n7), .C(n30734), .D(n29574), 
         .Z(n2747)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_226.init = 16'h0020;
    LUT4 Select_4291_i2_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31466), 
         .C(\read_value[6]_adj_77 ), .D(n33385), .Z(n2_adj_78)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4291_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_1554_i3_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[2]), 
         .D(n224[2]), .Z(n3922[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_440 (.A(sendcount[0]), .B(\sendcount[1] ), .Z(n31584)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i1_2_lut_rep_440.init = 16'h8888;
    LUT4 Select_4294_i2_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31466), 
         .C(\read_value[3]_adj_79 ), .D(rw), .Z(n2_adj_80)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4294_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_1554_i2_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[1]), 
         .D(n224[1]), .Z(n3922[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 i14821_3_lut_4_lut (.A(sendcount[0]), .B(\sendcount[1] ), .C(n9_adj_53), 
         .D(sendcount[2]), .Z(n17[2])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i14821_3_lut_4_lut.init = 16'h7f8f;
    LUT4 i14749_2_lut_rep_441 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n31585)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14749_2_lut_rep_441.init = 16'heeee;
    LUT4 i2_2_lut (.A(esc_data[7]), .B(esc_data[0]), .Z(n7)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_2_lut.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_391_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(sendcount[2]), 
         .Z(n31535)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam i1_2_lut_rep_391_3_lut.init = 16'h1e1e;
    LUT4 i3396_2_lut_rep_442 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n31586)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i3396_2_lut_rep_442.init = 16'h9999;
    LUT4 Select_4295_i2_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31466), 
         .C(\read_value[2]_adj_81 ), .D(rw), .Z(n2_adj_82)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4295_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4297_i2_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(n31466), 
         .C(\read_value[0]_adj_83 ), .D(n33385), .Z(n2_adj_84)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_4297_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_522_i4_3_lut (.A(n2747), .B(esc_data[3]), .C(n1474[18]), 
         .Z(n2216[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_522_i4_3_lut.init = 16'hcaca;
    PFUMX i22642 (.BLUT(n30707), .ALUT(n13_adj_151), .C0(n5834), .Z(n30708));
    LUT4 mux_522_i2_3_lut (.A(n2747), .B(esc_data[1]), .C(n1474[18]), 
         .Z(n2216[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_522_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1599_i1_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[0]), 
         .D(n224_adj_91[0]), .Z(n4095[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1599_i19_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[18]), 
         .D(n224_adj_91[18]), .Z(n4095[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 i14822_2_lut_2_lut_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(n9_adj_53), .Z(n17[1])) /* synthesis lut_function=(!(A (B (C))+!A !(B+!(C)))) */ ;
    defparam i14822_2_lut_2_lut_3_lut.init = 16'h6f6f;
    LUT4 n13158_bdd_4_lut_22664_4_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(\buffer[5] [0]), .D(\buffer[4] [0]), .Z(n30706)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam n13158_bdd_4_lut_22664_4_lut.init = 16'h6420;
    LUT4 mux_1599_i32_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[31]), 
         .D(n224_adj_91[31]), .Z(n4095[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i32_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_522_i1_3_lut (.A(n2747), .B(esc_data[0]), .C(n1474[18]), 
         .Z(n2216[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_522_i1_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_adj_227 (.A(n27445), .B(\control_reg[7] ), .C(n31601), 
         .Z(n34)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_adj_227.init = 16'h0808;
    LUT4 i3_4_lut (.A(register_addr[1]), .B(register_addr[2]), .C(n31539), 
         .D(n29256), .Z(n29257)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i3_4_lut.init = 16'h0200;
    LUT4 mux_1554_i21_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[20]), 
         .D(n224[20]), .Z(n3922[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1599_i18_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[17]), 
         .D(n224_adj_91[17]), .Z(n4095[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1599_i31_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[30]), 
         .D(n224_adj_91[30]), .Z(n4095[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i31_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1554_i27_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[26]), 
         .D(n224[26]), .Z(n3922[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i27_3_lut_4_lut.init = 16'hf780;
    LUT4 i4438_3_lut (.A(n1474[19]), .B(n1474[18]), .C(busy), .Z(n11203)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4438_3_lut.init = 16'hcece;
    LUT4 i3_3_lut_4_lut (.A(n31428), .B(n31576), .C(n31497), .D(n19332), 
         .Z(n9331)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i3_3_lut_4_lut.init = 16'h0080;
    LUT4 mux_1554_i26_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[25]), 
         .D(n224[25]), .Z(n3922[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i26_3_lut_4_lut.init = 16'hf780;
    FD1P3AX reg_addr_i0_i7 (.D(\buffer[1] [7]), .SP(n2806), .CK(debug_c_c), 
            .Q(register_addr_c[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i7.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i6 (.D(\buffer[1] [6]), .SP(n2806), .CK(debug_c_c), 
            .Q(register_addr_c[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i6.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i5 (.D(\buffer[1] [5]), .SP(n2806), .CK(debug_c_c), 
            .Q(register_addr[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i5.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i4 (.D(\buffer[1] [4]), .SP(n2806), .CK(debug_c_c), 
            .Q(register_addr[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i4.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i3 (.D(\buffer[1] [3]), .SP(n2806), .CK(debug_c_c), 
            .Q(register_addr[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i3.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i2 (.D(\buffer[1] [2]), .SP(n2806), .CK(debug_c_c), 
            .Q(register_addr[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i2.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i1 (.D(\buffer[1] [1]), .SP(n2806), .CK(debug_c_c), 
            .Q(register_addr[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i1.GSR = "ENABLED";
    LUT4 i5582_3_lut (.A(busy), .B(n1486), .C(n1474[19]), .Z(n12350)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5582_3_lut.init = 16'ha8a8;
    LUT4 i1_2_lut_adj_228 (.A(sendcount[0]), .B(sendcount[3]), .Z(n13_adj_151)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_228.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_446 (.A(register_addr[5]), .B(register_addr[4]), .Z(n31590)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_446.init = 16'heeee;
    LUT4 i12433_3_lut (.A(\register[0][5] ), .B(expansion5_c), .C(register_addr[1]), 
         .Z(n79)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i12433_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_229 (.A(register_addr[1]), .B(\register[1][5] ), .Z(n159)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_229.init = 16'h4444;
    LUT4 i1_2_lut_adj_230 (.A(n1474[6]), .B(n1474[11]), .Z(n1927)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_230.init = 16'heeee;
    LUT4 i5_4_lut (.A(n9_adj_122), .B(n1474[15]), .C(n8), .D(n1474[1]), 
         .Z(debug_c_2)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_adj_231 (.A(n1489), .B(n1474[9]), .Z(n8)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_2_lut_adj_231.init = 16'heeee;
    LUT4 i1_4_lut_adj_232 (.A(n31549), .B(n1474[7]), .C(n10_adj_157), 
         .D(n31550), .Z(debug_c_3)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_232.init = 16'hfffe;
    LUT4 reduce_or_2659_i1_2_lut_3_lut_4_lut_4_lut (.A(n31478), .B(register_addr[0]), 
         .C(n31477), .D(register_addr[1]), .Z(n9379)) /* synthesis lut_function=(!(A ((C+(D))+!B))) */ ;
    defparam reduce_or_2659_i1_2_lut_3_lut_4_lut_4_lut.init = 16'h555d;
    LUT4 i1_2_lut_rep_362_3_lut_4_lut (.A(register_addr[5]), .B(register_addr[4]), 
         .C(n31596), .D(register_addr[3]), .Z(n31506)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_362_3_lut_4_lut.init = 16'hfffe;
    LUT4 i4_4_lut (.A(n1474[2]), .B(n1474[10]), .C(n1474[18]), .D(n1474[6]), 
         .Z(n10_adj_157)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 i3_4_lut_adj_233 (.A(\buffer[0] [3]), .B(\buffer[0] [5]), .C(\buffer[0] [4]), 
         .D(\buffer[0] [6]), .Z(n28917)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i3_4_lut_adj_233.init = 16'hfffe;
    LUT4 i1_2_lut_rep_272_3_lut_4_lut (.A(\select[4] ), .B(n31470), .C(n29492), 
         .D(prev_select_adj_85), .Z(n31416)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_272_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_adj_234 (.A(register_addr[1]), .B(\steps_reg[7] ), .Z(n11)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_234.init = 16'h8888;
    LUT4 i4_4_lut_adj_235 (.A(n1474[4]), .B(n31513), .C(n1486), .D(n6), 
         .Z(debug_c_4)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut_adj_235.init = 16'hfffe;
    LUT4 mux_1599_i17_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[16]), 
         .D(n224_adj_91[16]), .Z(n4095[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1599_i6_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[5]), 
         .D(n224_adj_91[5]), .Z(n4095[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1599_i16_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[15]), 
         .D(n224_adj_91[15]), .Z(n4095[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 i22014_2_lut_rep_452 (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .Z(n31596)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22014_2_lut_rep_452.init = 16'heeee;
    LUT4 i21908_2_lut_rep_400_3_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[5]), .Z(n31544)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i21908_2_lut_rep_400_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_371_3_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[4]), .Z(n31515)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_371_3_lut.init = 16'h1010;
    LUT4 i22075_3_lut_rep_380_4_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[4]), .D(register_addr[5]), .Z(n31524)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22075_3_lut_rep_380_4_lut.init = 16'hfffe;
    FD1P3IX buffer_0___i2 (.D(n28667), .SP(n13042), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i2.GSR = "ENABLED";
    FD1P3IX buffer_0___i3 (.D(n28659), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i3.GSR = "ENABLED";
    FD1P3IX buffer_0___i4 (.D(n28617), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i4.GSR = "ENABLED";
    FD1P3IX buffer_0___i5 (.D(n28615), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[0] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i5.GSR = "ENABLED";
    FD1P3IX buffer_0___i6 (.D(n28619), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[0] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i6.GSR = "ENABLED";
    FD1P3IX buffer_0___i7 (.D(n28621), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i7.GSR = "ENABLED";
    FD1P3IX buffer_0___i8 (.D(n28663), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i8.GSR = "ENABLED";
    FD1P3IX buffer_0___i9 (.D(n28613), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i9.GSR = "ENABLED";
    FD1P3IX buffer_0___i10 (.D(n28661), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i10.GSR = "ENABLED";
    FD1P3IX buffer_0___i11 (.D(n28625), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i11.GSR = "ENABLED";
    FD1P3IX buffer_0___i12 (.D(n28609), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i12.GSR = "ENABLED";
    FD1P3IX buffer_0___i13 (.D(n28611), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i13.GSR = "ENABLED";
    FD1P3IX buffer_0___i14 (.D(n28587), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i14.GSR = "ENABLED";
    FD1P3IX buffer_0___i15 (.D(n28623), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i15.GSR = "ENABLED";
    FD1P3IX buffer_0___i16 (.D(n28607), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i16.GSR = "ENABLED";
    FD1P3IX buffer_0___i17 (.D(n27602), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i17.GSR = "ENABLED";
    FD1P3IX buffer_0___i18 (.D(n27600), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i18.GSR = "ENABLED";
    FD1P3IX buffer_0___i19 (.D(n27603), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i19.GSR = "ENABLED";
    FD1P3IX buffer_0___i20 (.D(n27598), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[2] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i20.GSR = "ENABLED";
    FD1P3IX buffer_0___i21 (.D(n27539), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[2] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i21.GSR = "ENABLED";
    FD1P3IX buffer_0___i22 (.D(n27549), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[2] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i22.GSR = "ENABLED";
    FD1P3IX buffer_0___i23 (.D(n27557), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[2] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i23.GSR = "ENABLED";
    FD1P3IX buffer_0___i24 (.D(n27525), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[2] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i24.GSR = "ENABLED";
    FD1P3IX buffer_0___i25 (.D(n27505), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[3] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i25.GSR = "ENABLED";
    FD1P3IX buffer_0___i26 (.D(n27473), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[3] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i26.GSR = "ENABLED";
    FD1P3IX buffer_0___i27 (.D(n27533), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[3] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i27.GSR = "ENABLED";
    FD1P3IX buffer_0___i28 (.D(n27558), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[3] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i28.GSR = "ENABLED";
    FD1P3IX buffer_0___i29 (.D(n27492), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[3] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i29.GSR = "ENABLED";
    FD1P3IX buffer_0___i30 (.D(n27556), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[3] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i30.GSR = "ENABLED";
    FD1P3IX buffer_0___i31 (.D(n27555), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[3] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i31.GSR = "ENABLED";
    FD1P3IX buffer_0___i32 (.D(n27552), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[3] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i32.GSR = "ENABLED";
    FD1P3IX buffer_0___i33 (.D(n27551), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[4] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i33.GSR = "ENABLED";
    FD1P3IX buffer_0___i34 (.D(n27501), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[4] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i34.GSR = "ENABLED";
    FD1P3IX buffer_0___i35 (.D(n27544), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[4] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i35.GSR = "ENABLED";
    FD1P3IX buffer_0___i36 (.D(n27534), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[4] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i36.GSR = "ENABLED";
    FD1P3IX buffer_0___i37 (.D(n27427), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[4] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i37.GSR = "ENABLED";
    FD1P3IX buffer_0___i38 (.D(n27479), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[4] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i38.GSR = "ENABLED";
    FD1P3IX buffer_0___i39 (.D(n27611), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[4] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i39.GSR = "ENABLED";
    FD1P3IX buffer_0___i40 (.D(n27497), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[4] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i40.GSR = "ENABLED";
    FD1P3IX buffer_0___i41 (.D(n27514), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[5] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i41.GSR = "ENABLED";
    FD1P3IX buffer_0___i42 (.D(n27513), .SP(n9472), .CD(n31473), .CK(debug_c_c), 
            .Q(\buffer[5] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i42.GSR = "ENABLED";
    FD1P3IX buffer_0___i43 (.D(n27477), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[5] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i43.GSR = "ENABLED";
    FD1P3IX buffer_0___i44 (.D(n27512), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[5] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i44.GSR = "ENABLED";
    FD1P3IX buffer_0___i45 (.D(n27511), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[5] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i45.GSR = "ENABLED";
    FD1P3IX buffer_0___i46 (.D(n27466), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[5] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i46.GSR = "ENABLED";
    FD1P3IX buffer_0___i47 (.D(n27506), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[5] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i47.GSR = "ENABLED";
    FD1P3IX buffer_0___i48 (.D(n27500), .SP(n9472), .CD(n33390), .CK(debug_c_c), 
            .Q(\buffer[5] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i48.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_389_3_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[5]), .Z(n31533)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_389_3_lut.init = 16'hfefe;
    LUT4 i4385_2_lut_rep_358_3_lut_4_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[4]), .D(register_addr[5]), .Z(n31502)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i4385_2_lut_rep_358_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_395_3_lut (.A(register_addr_c[7]), .B(register_addr_c[6]), 
         .C(register_addr[3]), .Z(n31539)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_395_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_236 (.A(n45_adj_163), .B(n112), .C(register_addr[0]), 
         .D(n28900), .Z(n6006)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B))) */ ;
    defparam i1_4_lut_adj_236.init = 16'h333b;
    LUT4 i1_2_lut_3_lut_adj_237 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n29361)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_237.init = 16'hfbfb;
    LUT4 i18001_3_lut (.A(n31601), .B(\register[2] [0]), .C(register_addr[1]), 
         .Z(n45_adj_163)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i18001_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_238 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n29362)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_238.init = 16'hbfbf;
    LUT4 i4_4_lut_adj_239 (.A(n1474[11]), .B(n1474[8]), .C(n1474[13]), 
         .D(n1474[10]), .Z(n10)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut_adj_239.init = 16'hfffe;
    LUT4 i1_2_lut_adj_240 (.A(register_addr[1]), .B(\steps_reg[5] ), .Z(n14_adj_86)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_240.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_241 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n29358)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_241.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_242 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n29359)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_242.init = 16'hbfbf;
    LUT4 mux_1599_i15_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[14]), 
         .D(n224_adj_91[14]), .Z(n4095[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1599_i14_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[13]), 
         .D(n224_adj_91[13]), .Z(n4095[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i37_3_lut (.A(\register[0][4] ), .B(expansion4_out), .C(register_addr[1]), 
         .Z(n25)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i37_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_456 (.A(n1474[3]), .B(debug_c_7), .Z(n31600)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_456.init = 16'h8888;
    LUT4 i1_2_lut_adj_243 (.A(register_addr[1]), .B(\register[1][4] ), .Z(n19)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_2_lut_adj_243.init = 16'h4444;
    LUT4 mux_1599_i5_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[4]), 
         .D(n224_adj_91[4]), .Z(n4095[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_3_lut_rep_457 (.A(force_pause), .B(\register[0][2] ), .C(timeout_pause), 
         .Z(n31601)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[6:17])
    defparam i2_3_lut_rep_457.init = 16'hfefe;
    LUT4 mux_1599_i4_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[3]), 
         .D(n224_adj_91[3]), .Z(n4095[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1599_i3_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[2]), 
         .D(n224_adj_91[2]), .Z(n4095[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_244 (.A(register_addr[1]), .B(\steps_reg[6] ), .Z(n13_adj_87)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_244.init = 16'h8888;
    LUT4 i15238_2_lut_rep_393_4_lut (.A(force_pause), .B(\register[0][2] ), 
         .C(timeout_pause), .D(\register[0][7] ), .Z(n31537)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[6:17])
    defparam i15238_2_lut_rep_393_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_4_lut_adj_245 (.A(force_pause), .B(\register[0][2] ), 
         .C(timeout_pause), .D(clk_1Hz), .Z(signal_light_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[6:17])
    defparam i1_2_lut_4_lut_adj_245.init = 16'hfffe;
    LUT4 i22319_2_lut_2_lut (.A(n31501), .B(n13042), .Z(n9472)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i22319_2_lut_2_lut.init = 16'hdddd;
    LUT4 mux_1599_i2_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[1]), 
         .D(n224_adj_91[1]), .Z(n4095[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_246 (.A(register_addr[1]), .B(\steps_reg[3] ), .Z(n12)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_246.init = 16'h8888;
    LUT4 i22_3_lut (.A(\control_reg[4] ), .B(\div_factor_reg[4] ), .C(register_addr[1]), 
         .Z(n12_adj_172)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i22_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_247 (.A(register_addr[1]), .B(\steps_reg[4] ), .Z(n6_adj_173)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_2_lut_adj_247.init = 16'h8888;
    LUT4 i1_4_lut_adj_248 (.A(n29163), .B(debug_c_7), .C(n1474[0]), .D(n1474[1]), 
         .Z(n13789)) /* synthesis lut_function=(A+!(B+!(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_248.init = 16'hbbba;
    LUT4 i3_4_lut_adj_249 (.A(sendcount[3]), .B(n31585), .C(sendcount[2]), 
         .D(n31581), .Z(n29163)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_249.init = 16'h0200;
    LUT4 i1_2_lut_adj_250 (.A(register_addr[0]), .B(\control_reg[7]_adj_88 ), 
         .Z(n8636)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_250.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_251 (.A(n31571), .B(n31424), .C(register_addr[0]), 
         .D(n31512), .Z(n13948)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A (C+!(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_251.init = 16'h0f02;
    LUT4 i1_2_lut_3_lut_4_lut_adj_252 (.A(n31571), .B(n31424), .C(register_addr[0]), 
         .D(n31512), .Z(n12369)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_252.init = 16'hf020;
    LUT4 mux_1599_i13_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[12]), 
         .D(n224_adj_91[12]), .Z(n4095[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1554_i23_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[22]), 
         .D(n224[22]), .Z(n3922[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 i21940_2_lut (.A(n33385), .B(register_addr[5]), .Z(n29492)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21940_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_253 (.A(prev_select_adj_85), .B(n29170), .C(n29492), 
         .D(n31466), .Z(n9301)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i3_4_lut_adj_253.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_254 (.A(n31596), .B(n31507), .C(n31512), 
         .D(n29231), .Z(n14523)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_254.init = 16'hf1f0;
    FD1S3IX state_FSM_i2 (.D(n28693), .CK(debug_c_c), .CD(n33390), .Q(n1474[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i2.GSR = "ENABLED";
    LUT4 i2_3_lut_adj_255 (.A(n29231), .B(n35), .C(register_addr[4]), 
         .Z(n4007)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i2_3_lut_adj_255.init = 16'h0808;
    LUT4 n79_bdd_4_lut (.A(n79), .B(n159), .C(register_addr[0]), .D(n31487), 
         .Z(n31407)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n79_bdd_4_lut.init = 16'h00ca;
    LUT4 i2_4_lut_adj_256 (.A(n31479), .B(register_addr[5]), .C(\select[4] ), 
         .D(rw), .Z(n29231)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i2_4_lut_adj_256.init = 16'h0040;
    LUT4 mux_1599_i30_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[29]), 
         .D(n224_adj_91[29]), .Z(n4095[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i30_3_lut_4_lut.init = 16'hf780;
    FD1P3IX tx_data_i0_i2 (.D(esc_data[2]), .SP(n31469), .CD(n16770), 
            .CK(debug_c_c), .Q(tx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i5 (.D(esc_data[5]), .SP(n31469), .CD(n16770), 
            .CK(debug_c_c), .Q(tx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i6 (.D(esc_data[6]), .SP(n31469), .CD(n16770), 
            .CK(debug_c_c), .Q(tx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i7 (.D(esc_data[7]), .SP(n31469), .CD(n16770), 
            .CK(debug_c_c), .Q(tx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i3 (.D(n9241[3]), .SP(n13834), .CD(n16768), .CK(debug_c_c), 
            .Q(esc_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i3.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i5 (.D(n9241[5]), .SP(n13834), .CD(n16768), .CK(debug_c_c), 
            .Q(esc_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i5.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i6 (.D(n9241[6]), .SP(n13834), .CD(n16768), .CK(debug_c_c), 
            .Q(esc_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i6.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i7 (.D(n9241[7]), .SP(n13834), .CD(n16768), .CK(debug_c_c), 
            .Q(esc_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i7.GSR = "ENABLED";
    LUT4 i2_2_lut_4_lut_4_lut (.A(n31478), .B(n31477), .C(register_addr[0]), 
         .D(register_addr[1]), .Z(n27680)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D))))) */ ;
    defparam i2_2_lut_4_lut_4_lut.init = 16'h5775;
    LUT4 i2_3_lut_adj_257 (.A(n27484), .B(\control_reg[7]_adj_88 ), .C(n31601), 
         .Z(n32_adj_89)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_adj_257.init = 16'h0808;
    LUT4 i9993_2_lut_3_lut_4_lut_4_lut (.A(n31478), .B(n14454), .C(n31477), 
         .D(register_addr[1]), .Z(n16765)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B))) */ ;
    defparam i9993_2_lut_3_lut_4_lut_4_lut.init = 16'h4c44;
    FD1S3IX state_FSM_i3 (.D(n13465), .CK(debug_c_c), .CD(n33390), .Q(n1474[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i3.GSR = "ENABLED";
    FD1S3IX state_FSM_i4 (.D(n12482), .CK(debug_c_c), .CD(n33390), .Q(n1474[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i4.GSR = "ENABLED";
    FD1S3IX state_FSM_i5 (.D(n29229), .CK(debug_c_c), .CD(n33390), .Q(n1474[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i5.GSR = "ENABLED";
    FD1S3IX state_FSM_i6 (.D(n29205), .CK(debug_c_c), .CD(n33390), .Q(n1474[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i6.GSR = "ENABLED";
    FD1S3IX state_FSM_i7 (.D(n1474[5]), .CK(debug_c_c), .CD(n33390), .Q(n1474[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i7.GSR = "ENABLED";
    FD1S3IX state_FSM_i8 (.D(n1474[6]), .CK(debug_c_c), .CD(n33390), .Q(n1474[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i8.GSR = "ENABLED";
    FD1S3IX state_FSM_i9 (.D(n1474[7]), .CK(debug_c_c), .CD(n33390), .Q(n1474[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i9.GSR = "ENABLED";
    FD1S3IX state_FSM_i10 (.D(n1474[8]), .CK(debug_c_c), .CD(n33390), 
            .Q(n1474[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i10.GSR = "ENABLED";
    FD1S3IX state_FSM_i11 (.D(n1579), .CK(debug_c_c), .CD(n33390), .Q(n1474[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i11.GSR = "ENABLED";
    FD1S3IX state_FSM_i12 (.D(n1474[10]), .CK(debug_c_c), .CD(n33390), 
            .Q(n1474[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i12.GSR = "ENABLED";
    FD1S3IX state_FSM_i13 (.D(n1474[11]), .CK(debug_c_c), .CD(n33390), 
            .Q(n1474[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i13.GSR = "ENABLED";
    FD1S3IX state_FSM_i14 (.D(n1474[12]), .CK(debug_c_c), .CD(n33390), 
            .Q(n1474[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i14.GSR = "ENABLED";
    FD1S3IX state_FSM_i15 (.D(n1585), .CK(debug_c_c), .CD(n33390), .Q(n1492));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i15.GSR = "ENABLED";
    FD1S3IX state_FSM_i16 (.D(n1586), .CK(debug_c_c), .CD(n33390), .Q(n1474[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i16.GSR = "ENABLED";
    FD1S3IX state_FSM_i17 (.D(n11217), .CK(debug_c_c), .CD(n33390), .Q(n1474[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i17.GSR = "ENABLED";
    FD1S3IX state_FSM_i18 (.D(n12348), .CK(debug_c_c), .CD(n33390), .Q(n1489));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i18.GSR = "ENABLED";
    FD1S3IX state_FSM_i19 (.D(n28605), .CK(debug_c_c), .CD(n33390), .Q(n1474[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i19.GSR = "ENABLED";
    FD1S3IX state_FSM_i20 (.D(n11203), .CK(debug_c_c), .CD(n33390), .Q(n1474[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i20.GSR = "ENABLED";
    FD1S3IX state_FSM_i21 (.D(n12350), .CK(debug_c_c), .CD(n33390), .Q(n1486));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i21.GSR = "ENABLED";
    LUT4 mux_1599_i29_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[28]), 
         .D(n224_adj_91[28]), .Z(n4095[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i29_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1599_i28_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[27]), 
         .D(n224_adj_91[27]), .Z(n4095[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i28_3_lut_4_lut.init = 16'hf780;
    FD1P3AX rw_498_rep_466 (.D(n1474[10]), .SP(n2806), .CK(debug_c_c), 
            .Q(n33385));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498_rep_466.GSR = "ENABLED";
    LUT4 mux_1599_i27_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[26]), 
         .D(n224_adj_91[26]), .Z(n4095[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i27_3_lut_4_lut.init = 16'hf780;
    LUT4 i5_4_lut_adj_258 (.A(n9), .B(\select[4] ), .C(n8_adj_182), .D(register_addr[4]), 
         .Z(n9305)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i5_4_lut_adj_258.init = 16'h0080;
    LUT4 mux_1599_i26_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[25]), 
         .D(n224_adj_91[25]), .Z(n4095[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i26_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_2_lut_adj_259 (.A(register_addr[5]), .B(prev_select_adj_6), 
         .Z(n8_adj_182)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_2_lut_adj_259.init = 16'h2222;
    LUT4 i15043_3_lut_4_lut (.A(n31476), .B(n1492), .C(n9_adj_53), .D(sendcount[0]), 
         .Z(n15[0])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (C (D)))) */ ;
    defparam i15043_3_lut_4_lut.init = 16'h0ddd;
    LUT4 i1_2_lut_adj_260 (.A(register_addr[5]), .B(register_addr[4]), .Z(n29256)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_260.init = 16'h8888;
    LUT4 i2_3_lut_rep_283_4_lut (.A(register_addr[1]), .B(n31477), .C(n31465), 
         .D(prev_select_adj_90), .Z(n31427)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_283_4_lut.init = 16'h00e0;
    LUT4 i1_2_lut_adj_261 (.A(register_addr[0]), .B(register_addr[1]), .Z(n19332)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_261.init = 16'hbbbb;
    LUT4 mux_1599_i25_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[24]), 
         .D(n224_adj_91[24]), .Z(n4095[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i25_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_262 (.A(n31523), .B(debug_c_7), .C(n13490), .D(n8_adj_185), 
         .Z(n28693)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_262.init = 16'hdc50;
    LUT4 i1_3_lut (.A(n31454), .B(n1474[1]), .C(n1474[0]), .Z(n8_adj_185)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut.init = 16'hecec;
    LUT4 i4_4_lut_adj_263 (.A(n7_adj_186), .B(n29277), .C(rx_data[2]), 
         .D(rx_data[0]), .Z(n13490)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i4_4_lut_adj_263.init = 16'h8000;
    LUT4 i9992_2_lut_3_lut_4_lut_4_lut (.A(n31478), .B(n14454), .C(n31477), 
         .D(register_addr[1]), .Z(n16764)) /* synthesis lut_function=(A (B (C+!(D)))) */ ;
    defparam i9992_2_lut_3_lut_4_lut_4_lut.init = 16'h8088;
    LUT4 i2_4_lut_adj_264 (.A(escape), .B(n31600), .C(n29648), .D(rx_data[6]), 
         .Z(n7_adj_186)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i2_4_lut_adj_264.init = 16'h0004;
    LUT4 i22089_3_lut (.A(rx_data[5]), .B(rx_data[7]), .C(rx_data[3]), 
         .Z(n29648)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22089_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_265 (.A(n1474[4]), .B(\buffer[0] [0]), .C(n11_c), 
         .D(n14_c), .Z(n28593)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_265.init = 16'heca0;
    LUT4 reduce_or_463_i1_3_lut_4_lut (.A(n31523), .B(n13490), .C(\buffer[0] [7]), 
         .D(n1474[9]), .Z(n1579)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(158[15] 160[18])
    defparam reduce_or_463_i1_3_lut_4_lut.init = 16'hff80;
    PFUMX i38 (.BLUT(n25), .ALUT(n19), .C0(register_addr[0]), .Z(n28));
    LUT4 i1_4_lut_adj_266 (.A(n5834), .B(n13_adj_151), .C(n31501), .D(n1492), 
         .Z(n16768)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_266.init = 16'h8000;
    LUT4 mux_429_Mux_3_i4_3_lut (.A(\buffer[4] [3]), .B(\buffer[5] [3]), 
         .C(sendcount[0]), .Z(n4_adj_57)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_3_i4_3_lut.init = 16'hacac;
    LUT4 esc_data_2__bdd_4_lut (.A(esc_data[2]), .B(esc_data[1]), .C(esc_data[3]), 
         .D(esc_data[4]), .Z(n30734)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C (D))+!B !(C+(D))))) */ ;
    defparam esc_data_2__bdd_4_lut.init = 16'h4801;
    LUT4 mux_429_Mux_5_i4_3_lut (.A(\buffer[4] [5]), .B(\buffer[5] [5]), 
         .C(sendcount[0]), .Z(n4_adj_56)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_5_i4_3_lut.init = 16'hacac;
    LUT4 mux_429_Mux_6_i4_3_lut (.A(\buffer[4] [6]), .B(\buffer[5] [6]), 
         .C(sendcount[0]), .Z(n4_adj_55)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_6_i4_3_lut.init = 16'hacac;
    LUT4 mux_429_Mux_7_i4_3_lut (.A(\buffer[4] [7]), .B(\buffer[5] [7]), 
         .C(sendcount[0]), .Z(n4_c)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_7_i4_3_lut.init = 16'hacac;
    LUT4 i1_4_lut_adj_267 (.A(\register[2] [3]), .B(n112), .C(n19332), 
         .D(n28900), .Z(n6003)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B))) */ ;
    defparam i1_4_lut_adj_267.init = 16'h333b;
    LUT4 i1_4_lut_adj_268 (.A(register_addr[1]), .B(n31506), .C(register_addr[0]), 
         .D(register_addr[2]), .Z(n112)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_4_lut_adj_268.init = 16'hfeff;
    LUT4 i2_3_lut_adj_269 (.A(register_addr[2]), .B(register_addr[3]), .C(n31524), 
         .Z(n28900)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_adj_269.init = 16'hfefe;
    LUT4 i22355_4_lut (.A(n31539), .B(n31590), .C(register_addr[2]), .D(n31591), 
         .Z(n27428)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;
    defparam i22355_4_lut.init = 16'h0111;
    LUT4 mux_1599_i24_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[23]), 
         .D(n224_adj_91[23]), .Z(n4095[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1554_i25_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[24]), 
         .D(n224[24]), .Z(n3922[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i25_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1554_i24_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[23]), 
         .D(n224[23]), .Z(n3922[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1599_i23_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[22]), 
         .D(n224_adj_91[22]), .Z(n4095[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1599_i22_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[21]), 
         .D(n224_adj_91[21]), .Z(n4095[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1554_i20_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[19]), 
         .D(n224[19]), .Z(n3922[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i20_3_lut_4_lut.init = 16'hf780;
    PFUMX i21 (.BLUT(n12_adj_172), .ALUT(n6_adj_173), .C0(register_addr[0]), 
          .Z(n28827));
    LUT4 i1_2_lut_adj_270 (.A(register_addr[0]), .B(\control_reg[7]_adj_37 ), 
         .Z(n8654)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_270.init = 16'h4444;
    LUT4 mux_1599_i21_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[20]), 
         .D(n224_adj_91[20]), .Z(n4095[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 i22323_4_lut (.A(n7_adj_125), .B(n29560), .C(n31552), .D(n1474[3]), 
         .Z(n13042)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C+!(D))))) */ ;
    defparam i22323_4_lut.init = 16'h0544;
    LUT4 i22006_3_lut (.A(n1474[13]), .B(n1474[0]), .C(n1474[4]), .Z(n29560)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22006_3_lut.init = 16'hfefe;
    LUT4 mux_1599_i12_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[11]), 
         .D(n224_adj_91[11]), .Z(n4095[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1599_i11_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[10]), 
         .D(n224_adj_91[10]), .Z(n4095[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1599_i10_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[9]), 
         .D(n224_adj_91[9]), .Z(n4095[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1599_i9_3_lut_4_lut (.A(n31416), .B(n31423), .C(databus[8]), 
         .D(n224_adj_91[8]), .Z(n4095[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1599_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1554_i22_3_lut_4_lut (.A(n31415), .B(n31423), .C(databus[21]), 
         .D(n224[21]), .Z(n3922[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1554_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_271 (.A(n29424), .B(n31600), .C(escape), .D(n30736), 
         .Z(n29229)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_271.init = 16'hccc8;
    LUT4 reduce_or_469_i1_3_lut (.A(busy), .B(n1474[13]), .C(n1486), .Z(n1585)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam reduce_or_469_i1_3_lut.init = 16'hdcdc;
    LUT4 i471_2_lut (.A(n5834), .B(n1492), .Z(n1586)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i471_2_lut.init = 16'h4444;
    PFUMX i23004 (.BLUT(n31645), .ALUT(n31646), .C0(n1927), .Z(n31647));
    PFUMX i23002 (.BLUT(n31642), .ALUT(n31643), .C0(n1927), .Z(n31644));
    PFUMX i23000 (.BLUT(n31639), .ALUT(n31640), .C0(sendcount[0]), .Z(n31641));
    PFUMX i22998 (.BLUT(n31636), .ALUT(n31637), .C0(sendcount[0]), .Z(n31638));
    PFUMX i22996 (.BLUT(n31633), .ALUT(n31634), .C0(sendcount[0]), .Z(n31635));
    PFUMX i22994 (.BLUT(n31630), .ALUT(n31631), .C0(sendcount[0]), .Z(n31632));
    PFUMX i22992 (.BLUT(n31627), .ALUT(n31628), .C0(sendcount[0]), .Z(n31629));
    PFUMX i22990 (.BLUT(n31624), .ALUT(n31625), .C0(sendcount[0]), .Z(n31626));
    LUT4 i1_2_lut_adj_272 (.A(rx_data[5]), .B(rx_data[0]), .Z(n29424)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_272.init = 16'hbbbb;
    PFUMX i22988 (.BLUT(n31621), .ALUT(n31622), .C0(sendcount[0]), .Z(n31623));
    LUT4 i4452_3_lut (.A(n1474[16]), .B(n2747), .C(busy), .Z(n11217)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4452_3_lut.init = 16'hcece;
    PFUMX i22986 (.BLUT(n31618), .ALUT(n31619), .C0(sendcount[3]), .Z(n5834));
    LUT4 i5581_3_lut (.A(busy), .B(n1489), .C(n1474[16]), .Z(n12348)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5581_3_lut.init = 16'ha8a8;
    LUT4 i2_4_lut_adj_273 (.A(n38), .B(busy), .C(n30342), .D(n1489), 
         .Z(n28605)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_273.init = 16'hfbfa;
    PFUMX i22982 (.BLUT(n31612), .ALUT(n31613), .C0(sendcount[0]), .Z(n31614));
    PFUMX i22980 (.BLUT(n31609), .ALUT(n31610), .C0(n31451), .Z(n31611));
    \UARTTransmitter(baud_div=12)  uart_output (.n33390(n33390), .tx_data({tx_data}), 
            .send(send), .\state[3] (\state[3] ), .\state[1] (\state[1] ), 
            .\state[0] (\state[0] ), .n1156(n1156), .n73(n73), .n31501(n31501), 
            .busy(busy), .n31473(n31473), .\reset_count[7] (\reset_count[7] ), 
            .\reset_count[6] (\reset_count[6] ), .\reset_count[5] (\reset_count[5] ), 
            .n27250(n27250), .uart_tx_c(uart_tx_c), .debug_c_c(debug_c_c), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(65[30] 70[52])
    \UARTReceiver(baud_div=12)  uart_input (.debug_c_c(debug_c_c), .n31501(n31501), 
            .rx_data({rx_data}), .n33390(n33390), .uart_rx_c(uart_rx_c), 
            .debug_c_7(debug_c_7), .n29424(n29424), .n29277(n29277), .n57(n57_adj_109), 
            .n31454(n31454), .n30736(n30736), .n31473(n31473), .n1502(n1474[4]), 
            .n1504(n1474[2]), .n13465(n13465), .n1506(n1474[0]), .escape(escape), 
            .n1503(n1474[3]), .n12482(n12482), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(60[27] 64[39])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=12) 
//

module \UARTTransmitter(baud_div=12)  (n33390, tx_data, send, \state[3] , 
            \state[1] , \state[0] , n1156, n73, n31501, busy, n31473, 
            \reset_count[7] , \reset_count[6] , \reset_count[5] , n27250, 
            uart_tx_c, debug_c_c, GND_net) /* synthesis syn_module_defined=1 */ ;
    input n33390;
    input [7:0]tx_data;
    input send;
    input \state[3] ;
    input \state[1] ;
    input \state[0] ;
    input n1156;
    output n73;
    input n31501;
    output busy;
    input n31473;
    input \reset_count[7] ;
    input \reset_count[6] ;
    input \reset_count[5] ;
    output n27250;
    output uart_tx_c;
    input debug_c_c;
    input GND_net;
    
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [3:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n30446, n30318;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n9451, n30770, n14987, n31188, n31598, n31187, n42, n29732, 
        n29733, n30317, n30316, n28969, n31315, n7, n10, n104, 
        n12, n28972, n40, n29734, n2;
    
    LUT4 state_1__bdd_4_lut_22674 (.A(state[1]), .B(state[0]), .C(state[3]), 
         .D(state[2]), .Z(n30446)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C (D))+!B (C (D)+!C !(D))))) */ ;
    defparam state_1__bdd_4_lut_22674.init = 16'h0f7e;
    FD1S3IX state__i0 (.D(n30318), .CK(bclk), .CD(n33390), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n9451), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    LUT4 state_1__bdd_4_lut (.A(state[1]), .B(state[3]), .C(state[0]), 
         .D(send), .Z(n30770)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+(C+(D))))) */ ;
    defparam state_1__bdd_4_lut.init = 16'h7ffe;
    LUT4 i71_4_lut_4_lut (.A(\state[3] ), .B(\state[1] ), .C(\state[0] ), 
         .D(n1156), .Z(n73)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;
    defparam i71_4_lut_4_lut.init = 16'h8001;
    LUT4 i1_2_lut_2_lut_3_lut (.A(n30770), .B(state[2]), .C(n31501), .Z(n14987)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_2_lut_3_lut.init = 16'hefef;
    FD1P3IX busy_34 (.D(n31598), .SP(n31188), .CD(n31473), .CK(bclk), 
            .Q(busy));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam busy_34.GSR = "ENABLED";
    LUT4 n31187_bdd_2_lut (.A(n31187), .B(state[2]), .Z(n31188)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n31187_bdd_2_lut.init = 16'h2222;
    LUT4 send_bdd_4_lut (.A(send), .B(state[0]), .C(state[1]), .D(state[3]), 
         .Z(n31187)) /* synthesis lut_function=(A (B (C (D))+!B !(C+(D)))+!A (B (C (D)))) */ ;
    defparam send_bdd_4_lut.init = 16'hc002;
    LUT4 i1_2_lut (.A(state[1]), .B(state[0]), .Z(n42)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i22172_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n29732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22172_3_lut.init = 16'hcaca;
    LUT4 i22173_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n29733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22173_3_lut.init = 16'hcaca;
    LUT4 state_3__bdd_4_lut (.A(state[3]), .B(state[0]), .C(send), .D(state[1]), 
         .Z(n30317)) /* synthesis lut_function=(A ((C (D))+!B)+!A !(B+!(C+(D)))) */ ;
    defparam state_3__bdd_4_lut.init = 16'hb332;
    LUT4 state_3__bdd_2_lut (.A(state[3]), .B(state[0]), .Z(n30316)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_3__bdd_2_lut.init = 16'h1111;
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(state[0]), .C(n31501), .Z(n28969)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 n2802_bdd_4_lut (.A(n31501), .B(state[3]), .C(n42), .D(state[2]), 
         .Z(n31315)) /* synthesis lut_function=(!((B (D)+!B !(C (D)))+!A)) */ ;
    defparam n2802_bdd_4_lut.init = 16'h2088;
    LUT4 i2_3_lut (.A(\reset_count[7] ), .B(\reset_count[6] ), .C(\reset_count[5] ), 
         .Z(n27250)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    PFUMX Mux_22_i15 (.BLUT(n7), .ALUT(n10), .C0(state[3]), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;
    FD1P3AX state__i3 (.D(n31315), .SP(n14987), .CK(bclk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n9451), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n9451), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n9451), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n9451), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n9451), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n9451), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n9451), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    LUT4 i13088_1_lut_rep_454 (.A(state[3]), .Z(n31598)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i13088_1_lut_rep_454.init = 16'h5555;
    LUT4 i1_4_lut (.A(n31501), .B(state[3]), .C(n12), .D(state[2]), 
         .Z(n28972)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C))+!A)) */ ;
    defparam i1_4_lut.init = 16'h20a0;
    LUT4 i22_2_lut (.A(state[1]), .B(state[0]), .Z(n12)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i22_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_4_lut (.A(state[3]), .B(state[2]), .C(n42), .D(n31501), 
         .Z(n40)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i1_4_lut_4_lut.init = 16'h3400;
    PFUMX i22174 (.BLUT(n29732), .ALUT(n29733), .C0(state[1]), .Z(n29734));
    LUT4 Mux_22_i7_4_lut (.A(n2), .B(n29734), .C(state[2]), .D(state[1]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i15244_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i15244_4_lut.init = 16'hfcee;
    FD1P3AX state__i2 (.D(n40), .SP(n14987), .CK(bclk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    FD1P3AX state__i1 (.D(n28972), .SP(n14987), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    FD1P3JX tx_35 (.D(n104), .SP(n30446), .PD(n33390), .CK(bclk), .Q(uart_tx_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    LUT4 i3_4_lut (.A(send), .B(state[3]), .C(state[1]), .D(n28969), 
         .Z(n9451)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i3_4_lut.init = 16'h0200;
    PFUMX i22575 (.BLUT(n30317), .ALUT(n30316), .C0(state[2]), .Z(n30318));
    \ClockDividerP(factor=12)  baud_gen (.bclk(bclk), .debug_c_c(debug_c_c), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12) 
//

module \ClockDividerP(factor=12)  (bclk, debug_c_c, GND_net) /* synthesis syn_module_defined=1 */ ;
    output bclk;
    input debug_c_c;
    input GND_net;
    
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n8472, n27083, n27082;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n27081, n27080, n27079, n27078, n27077, n27076, n27075, 
        n27074, n27073, n27072, n27071, n27070, n27069, n27068, 
        n55, n56, n4, n16804, n52, n44, n35, n54, n48, n36, 
        n46, n32;
    wire [31:0]n102;
    
    wire n50, n40, n27019, n27018, n27017, n27016, n27015, n27014, 
        n27013, n27012, n27011, n27010, n27009, n27008, n27007, 
        n27006, n27005, n27004;
    
    FD1S3AX clk_o_14 (.D(n8472), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D sub_2086_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27083), .S0(n8472));
    defparam sub_2086_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2086_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2086_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2086_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27082), .COUT(n27083));
    defparam sub_2086_add_2_32.INIT0 = 16'h5555;
    defparam sub_2086_add_2_32.INIT1 = 16'h5555;
    defparam sub_2086_add_2_32.INJECT1_0 = "NO";
    defparam sub_2086_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27081), .COUT(n27082));
    defparam sub_2086_add_2_30.INIT0 = 16'h5555;
    defparam sub_2086_add_2_30.INIT1 = 16'h5555;
    defparam sub_2086_add_2_30.INJECT1_0 = "NO";
    defparam sub_2086_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27080), .COUT(n27081));
    defparam sub_2086_add_2_28.INIT0 = 16'h5555;
    defparam sub_2086_add_2_28.INIT1 = 16'h5555;
    defparam sub_2086_add_2_28.INJECT1_0 = "NO";
    defparam sub_2086_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27079), .COUT(n27080));
    defparam sub_2086_add_2_26.INIT0 = 16'h5555;
    defparam sub_2086_add_2_26.INIT1 = 16'h5555;
    defparam sub_2086_add_2_26.INJECT1_0 = "NO";
    defparam sub_2086_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27078), .COUT(n27079));
    defparam sub_2086_add_2_24.INIT0 = 16'h5555;
    defparam sub_2086_add_2_24.INIT1 = 16'h5555;
    defparam sub_2086_add_2_24.INJECT1_0 = "NO";
    defparam sub_2086_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27077), .COUT(n27078));
    defparam sub_2086_add_2_22.INIT0 = 16'h5555;
    defparam sub_2086_add_2_22.INIT1 = 16'h5555;
    defparam sub_2086_add_2_22.INJECT1_0 = "NO";
    defparam sub_2086_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27076), .COUT(n27077));
    defparam sub_2086_add_2_20.INIT0 = 16'h5555;
    defparam sub_2086_add_2_20.INIT1 = 16'h5555;
    defparam sub_2086_add_2_20.INJECT1_0 = "NO";
    defparam sub_2086_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27075), .COUT(n27076));
    defparam sub_2086_add_2_18.INIT0 = 16'h5555;
    defparam sub_2086_add_2_18.INIT1 = 16'h5555;
    defparam sub_2086_add_2_18.INJECT1_0 = "NO";
    defparam sub_2086_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27074), .COUT(n27075));
    defparam sub_2086_add_2_16.INIT0 = 16'h5555;
    defparam sub_2086_add_2_16.INIT1 = 16'h5555;
    defparam sub_2086_add_2_16.INJECT1_0 = "NO";
    defparam sub_2086_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27073), .COUT(n27074));
    defparam sub_2086_add_2_14.INIT0 = 16'h5555;
    defparam sub_2086_add_2_14.INIT1 = 16'h5555;
    defparam sub_2086_add_2_14.INJECT1_0 = "NO";
    defparam sub_2086_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27072), .COUT(n27073));
    defparam sub_2086_add_2_12.INIT0 = 16'h5555;
    defparam sub_2086_add_2_12.INIT1 = 16'h5555;
    defparam sub_2086_add_2_12.INJECT1_0 = "NO";
    defparam sub_2086_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27071), .COUT(n27072));
    defparam sub_2086_add_2_10.INIT0 = 16'h5555;
    defparam sub_2086_add_2_10.INIT1 = 16'h5555;
    defparam sub_2086_add_2_10.INJECT1_0 = "NO";
    defparam sub_2086_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27070), .COUT(n27071));
    defparam sub_2086_add_2_8.INIT0 = 16'h5555;
    defparam sub_2086_add_2_8.INIT1 = 16'h5555;
    defparam sub_2086_add_2_8.INJECT1_0 = "NO";
    defparam sub_2086_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27069), .COUT(n27070));
    defparam sub_2086_add_2_6.INIT0 = 16'h5555;
    defparam sub_2086_add_2_6.INIT1 = 16'h5555;
    defparam sub_2086_add_2_6.INJECT1_0 = "NO";
    defparam sub_2086_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27068), .COUT(n27069));
    defparam sub_2086_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2086_add_2_4.INIT1 = 16'h5555;
    defparam sub_2086_add_2_4.INJECT1_0 = "NO";
    defparam sub_2086_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_2086_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27068));
    defparam sub_2086_add_2_2.INIT0 = 16'h0000;
    defparam sub_2086_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2086_add_2_2.INJECT1_0 = "NO";
    defparam sub_2086_add_2_2.INJECT1_1 = "NO";
    LUT4 i22383_4_lut (.A(n55), .B(count[1]), .C(n56), .D(n4), .Z(n16804)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i22383_4_lut.init = 16'h0400;
    LUT4 i26_4_lut (.A(count[14]), .B(n52), .C(n44), .D(count[6]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i27_4_lut (.A(n35), .B(n54), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(count[3]), .B(count[0]), .Z(n4)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i23_4_lut (.A(count[24]), .B(n46), .C(n32), .D(count[16]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i15_3_lut (.A(count[15]), .B(count[31]), .C(count[5]), .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i17_4_lut (.A(count[26]), .B(count[12]), .C(count[28]), .D(count[18]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[13]), .B(count[22]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(count[20]), .B(count[4]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i6_2_lut.init = 16'heeee;
    FD1S3IX count_2679__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i0.GSR = "ENABLED";
    LUT4 i25_4_lut (.A(count[25]), .B(n50), .C(n40), .D(count[9]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(count[7]), .B(count[19]), .C(count[11]), .D(count[21]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[8]), .B(count[29]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i21_4_lut (.A(count[2]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i11_2_lut (.A(count[10]), .B(count[17]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i11_2_lut.init = 16'heeee;
    FD1S3IX count_2679__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i1.GSR = "ENABLED";
    FD1S3IX count_2679__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i2.GSR = "ENABLED";
    FD1S3IX count_2679__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i3.GSR = "ENABLED";
    FD1S3IX count_2679__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i4.GSR = "ENABLED";
    FD1S3IX count_2679__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i5.GSR = "ENABLED";
    FD1S3IX count_2679__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i6.GSR = "ENABLED";
    FD1S3IX count_2679__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i7.GSR = "ENABLED";
    FD1S3IX count_2679__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i8.GSR = "ENABLED";
    FD1S3IX count_2679__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i9.GSR = "ENABLED";
    FD1S3IX count_2679__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i10.GSR = "ENABLED";
    FD1S3IX count_2679__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i11.GSR = "ENABLED";
    FD1S3IX count_2679__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i12.GSR = "ENABLED";
    FD1S3IX count_2679__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i13.GSR = "ENABLED";
    FD1S3IX count_2679__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i14.GSR = "ENABLED";
    FD1S3IX count_2679__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i15.GSR = "ENABLED";
    FD1S3IX count_2679__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i16.GSR = "ENABLED";
    FD1S3IX count_2679__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i17.GSR = "ENABLED";
    FD1S3IX count_2679__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i18.GSR = "ENABLED";
    FD1S3IX count_2679__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i19.GSR = "ENABLED";
    FD1S3IX count_2679__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i20.GSR = "ENABLED";
    FD1S3IX count_2679__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i21.GSR = "ENABLED";
    FD1S3IX count_2679__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i22.GSR = "ENABLED";
    FD1S3IX count_2679__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i23.GSR = "ENABLED";
    FD1S3IX count_2679__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i24.GSR = "ENABLED";
    FD1S3IX count_2679__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i25.GSR = "ENABLED";
    FD1S3IX count_2679__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i26.GSR = "ENABLED";
    FD1S3IX count_2679__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i27.GSR = "ENABLED";
    FD1S3IX count_2679__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i28.GSR = "ENABLED";
    FD1S3IX count_2679__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i29.GSR = "ENABLED";
    FD1S3IX count_2679__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i30.GSR = "ENABLED";
    FD1S3IX count_2679__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n16804), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679__i31.GSR = "ENABLED";
    CCU2D count_2679_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27019), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_33.INIT1 = 16'h0000;
    defparam count_2679_add_4_33.INJECT1_0 = "NO";
    defparam count_2679_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27018), .COUT(n27019), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_31.INJECT1_0 = "NO";
    defparam count_2679_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27017), .COUT(n27018), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_29.INJECT1_0 = "NO";
    defparam count_2679_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27016), .COUT(n27017), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_27.INJECT1_0 = "NO";
    defparam count_2679_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27015), .COUT(n27016), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_25.INJECT1_0 = "NO";
    defparam count_2679_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27014), .COUT(n27015), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_23.INJECT1_0 = "NO";
    defparam count_2679_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27013), .COUT(n27014), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_21.INJECT1_0 = "NO";
    defparam count_2679_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27012), .COUT(n27013), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_19.INJECT1_0 = "NO";
    defparam count_2679_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27011), .COUT(n27012), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_17.INJECT1_0 = "NO";
    defparam count_2679_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27010), .COUT(n27011), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_15.INJECT1_0 = "NO";
    defparam count_2679_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27009), .COUT(n27010), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_13.INJECT1_0 = "NO";
    defparam count_2679_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27008), .COUT(n27009), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_11.INJECT1_0 = "NO";
    defparam count_2679_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27007), .COUT(n27008), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_9.INJECT1_0 = "NO";
    defparam count_2679_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27006), .COUT(n27007), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_7.INJECT1_0 = "NO";
    defparam count_2679_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27005), .COUT(n27006), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_5.INJECT1_0 = "NO";
    defparam count_2679_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27004), .COUT(n27005), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2679_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2679_add_4_3.INJECT1_0 = "NO";
    defparam count_2679_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2679_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27004), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2679_add_4_1.INIT0 = 16'hF000;
    defparam count_2679_add_4_1.INIT1 = 16'h0555;
    defparam count_2679_add_4_1.INJECT1_0 = "NO";
    defparam count_2679_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \UARTReceiver(baud_div=12) 
//

module \UARTReceiver(baud_div=12)  (debug_c_c, n31501, rx_data, n33390, 
            uart_rx_c, debug_c_7, n29424, n29277, n57, n31454, n30736, 
            n31473, n1502, n1504, n13465, n1506, escape, n1503, 
            n12482, GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n31501;
    output [7:0]rx_data;
    input n33390;
    input uart_rx_c;
    output debug_c_7;
    input n29424;
    input n29277;
    output n57;
    output n31454;
    output n30736;
    input n31473;
    input n1502;
    input n1504;
    output n13465;
    input n1506;
    input escape;
    input n1503;
    output n12482;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [7:0]rdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(22[12:17])
    
    wire n9399, n9401;
    wire [5:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    
    wire n28513, baud_reset, n19, n31561, n31520, n31498, n31491, 
        n31569, n31563, n13569, n19_adj_32, n30710, n30709, n31404;
    wire [7:0]n78;
    
    wire n13560, n13, n9415, n31603, n9417, n31568, n29323, n9419, 
        n9421, n29384, n9423, n22201, n9425, n9427, n10239, bclk, 
        n29203, n16637, n30789, n9429, n9431, n9433, n9435, n9437, 
        n9439, n29372, n24509, n19_adj_33, n9441, n27, n28297, 
        n31514, n29393, n31519, n30735, n31567, n31499, n25, n27_adj_34, 
        n28399, n21, n23, n28051, n16638, n4, n4_adj_35, n51, 
        n47;
    
    FD1P3AX rdata_i0_i0 (.D(n9399), .SP(n31501), .CK(debug_c_c), .Q(rdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i0.GSR = "ENABLED";
    FD1P3AX data_i0_i0 (.D(n9401), .SP(n31501), .CK(debug_c_c), .Q(rx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i0.GSR = "ENABLED";
    FD1S3IX state__i0 (.D(n28513), .CK(debug_c_c), .CD(n33390), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i0.GSR = "ENABLED";
    FD1S3JX baud_reset_52 (.D(n19), .CK(debug_c_c), .PD(n33390), .Q(baud_reset)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam baud_reset_52.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_354_4_lut (.A(state[4]), .B(state[3]), .C(n31561), 
         .D(n31520), .Z(n31498)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_354_4_lut.init = 16'heaff;
    LUT4 i1_2_lut_rep_347_4_lut (.A(state[4]), .B(state[3]), .C(n31561), 
         .D(state[5]), .Z(n31491)) /* synthesis lut_function=(!(A (D)+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_347_4_lut.init = 16'h00ea;
    LUT4 i2_3_lut_4_lut (.A(n31569), .B(n31563), .C(state[0]), .D(state[5]), 
         .Z(n13569)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i2_3_lut_4_lut.init = 16'h0100;
    LUT4 i2_3_lut_4_lut_adj_57 (.A(state[0]), .B(n31563), .C(state[5]), 
         .D(n31569), .Z(n19_adj_32)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_3_lut_4_lut_adj_57.init = 16'hffef;
    LUT4 n30710_bdd_4_lut (.A(n30710), .B(state[5]), .C(n30709), .D(state[0]), 
         .Z(n31404)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C (D))) */ ;
    defparam n30710_bdd_4_lut.init = 16'hf022;
    LUT4 i1_4_lut (.A(n78[1]), .B(rdata[1]), .C(n13560), .D(n13), .Z(n9415)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i4411_4_lut (.A(uart_rx_c), .B(rdata[1]), .C(n31569), .D(n31603), 
         .Z(n78[1])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4411_4_lut.init = 16'hcacc;
    LUT4 i1_4_lut_adj_58 (.A(n78[2]), .B(rdata[2]), .C(n13560), .D(n13), 
         .Z(n9417)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_58.init = 16'heca0;
    LUT4 i4409_4_lut (.A(uart_rx_c), .B(rdata[2]), .C(n31568), .D(n29323), 
         .Z(n78[2])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4409_4_lut.init = 16'hccca;
    LUT4 i1_2_lut (.A(state[3]), .B(state[2]), .Z(n29323)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_59 (.A(n78[3]), .B(rdata[3]), .C(n13560), .D(n13), 
         .Z(n9419)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_59.init = 16'heca0;
    LUT4 i4407_4_lut (.A(uart_rx_c), .B(rdata[3]), .C(n31603), .D(n29323), 
         .Z(n78[3])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4407_4_lut.init = 16'hccac;
    LUT4 i1_4_lut_adj_60 (.A(n78[4]), .B(rdata[4]), .C(n13560), .D(n13), 
         .Z(n9421)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_60.init = 16'heca0;
    LUT4 i4405_4_lut (.A(uart_rx_c), .B(rdata[4]), .C(state[2]), .D(n29384), 
         .Z(n78[4])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4405_4_lut.init = 16'hccca;
    LUT4 i1_4_lut_adj_61 (.A(n78[5]), .B(rdata[5]), .C(n13560), .D(n13), 
         .Z(n9423)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_61.init = 16'heca0;
    LUT4 i4403_4_lut (.A(uart_rx_c), .B(rdata[5]), .C(state[2]), .D(n22201), 
         .Z(n78[5])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4403_4_lut.init = 16'hcacc;
    LUT4 i1_4_lut_adj_62 (.A(n78[6]), .B(rdata[6]), .C(n13560), .D(n13), 
         .Z(n9425)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_62.init = 16'heca0;
    LUT4 i4401_4_lut (.A(uart_rx_c), .B(rdata[6]), .C(state[2]), .D(n29384), 
         .Z(n78[6])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4401_4_lut.init = 16'hccac;
    LUT4 i1_4_lut_adj_63 (.A(n78[7]), .B(rdata[7]), .C(n13560), .D(n13), 
         .Z(n9427)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_63.init = 16'heca0;
    LUT4 i1_4_lut_4_lut (.A(state[4]), .B(n10239), .C(bclk), .D(n31491), 
         .Z(n29203)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut.init = 16'h6a00;
    LUT4 i9865_3_lut_3_lut (.A(state[4]), .B(n10239), .C(bclk), .Z(n16637)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;
    defparam i9865_3_lut_3_lut.init = 16'ha6a6;
    LUT4 i4399_4_lut (.A(rdata[7]), .B(uart_rx_c), .C(state[2]), .D(n22201), 
         .Z(n78[7])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4399_4_lut.init = 16'hcaaa;
    LUT4 state_3__bdd_4_lut (.A(state[3]), .B(bclk), .C(state[2]), .D(state[1]), 
         .Z(n30789)) /* synthesis lut_function=(A (B+!(C (D)))+!A !(B+!(C (D)))) */ ;
    defparam state_3__bdd_4_lut.init = 16'h9aaa;
    LUT4 i1_4_lut_adj_64 (.A(rdata[1]), .B(rx_data[1]), .C(n13569), .D(n19_adj_32), 
         .Z(n9429)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_64.init = 16'heca0;
    LUT4 i1_4_lut_adj_65 (.A(rdata[2]), .B(rx_data[2]), .C(n13569), .D(n19_adj_32), 
         .Z(n9431)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_65.init = 16'heca0;
    LUT4 i1_4_lut_adj_66 (.A(rdata[3]), .B(rx_data[3]), .C(n13569), .D(n19_adj_32), 
         .Z(n9433)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_66.init = 16'heca0;
    LUT4 i1_4_lut_adj_67 (.A(rdata[4]), .B(rx_data[4]), .C(n13569), .D(n19_adj_32), 
         .Z(n9435)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_67.init = 16'heca0;
    LUT4 i1_4_lut_adj_68 (.A(rdata[5]), .B(rx_data[5]), .C(n13569), .D(n19_adj_32), 
         .Z(n9437)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_68.init = 16'heca0;
    LUT4 i1_4_lut_adj_69 (.A(rdata[6]), .B(rx_data[6]), .C(n13569), .D(n19_adj_32), 
         .Z(n9439)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_69.init = 16'heca0;
    LUT4 i22423_4_lut (.A(debug_c_7), .B(n29372), .C(uart_rx_c), .D(n24509), 
         .Z(n19_adj_33)) /* synthesis lut_function=(A (B+(C))+!A !((D)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i22423_4_lut.init = 16'ha8ec;
    LUT4 i1_4_lut_adj_70 (.A(rdata[7]), .B(rx_data[7]), .C(n13569), .D(n19_adj_32), 
         .Z(n9441)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_70.init = 16'heca0;
    LUT4 i43_4_lut (.A(state[5]), .B(n30789), .C(state[0]), .D(n27), 
         .Z(n28297)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i43_4_lut.init = 16'hc5c0;
    LUT4 i2_3_lut_4_lut_adj_71 (.A(n31514), .B(n29424), .C(rx_data[3]), 
         .D(n29277), .Z(n57)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_3_lut_4_lut_adj_71.init = 16'h1000;
    LUT4 i2_3_lut_rep_310_4_lut (.A(n31514), .B(n29424), .C(rx_data[1]), 
         .D(n29393), .Z(n31454)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_310_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut (.A(state[5]), .B(n31519), .C(state[0]), .D(bclk), 
         .Z(n28513)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_3_lut_4_lut.init = 16'hf400;
    LUT4 n30735_bdd_2_lut_3_lut (.A(rx_data[6]), .B(rx_data[7]), .C(n30735), 
         .Z(n30736)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam n30735_bdd_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_370_3_lut (.A(rx_data[6]), .B(rx_data[7]), .C(rx_data[2]), 
         .Z(n31514)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_370_3_lut.init = 16'hfefe;
    LUT4 i1_3_lut_4_lut_4_lut (.A(uart_rx_c), .B(n31520), .C(state[3]), 
         .D(n31519), .Z(n27)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A ((C (D))+!B)) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'hf131;
    FD1S3IX drdy_51 (.D(n19_adj_33), .CK(debug_c_c), .CD(n31473), .Q(debug_c_7));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam drdy_51.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_417 (.A(state[1]), .B(state[2]), .Z(n31561)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_rep_417.init = 16'h8888;
    LUT4 i1_3_lut_rep_375_4_lut (.A(state[1]), .B(state[2]), .C(state[3]), 
         .D(state[4]), .Z(n31519)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_3_lut_rep_375_4_lut.init = 16'hff80;
    LUT4 i1_2_lut_rep_419 (.A(state[1]), .B(state[4]), .Z(n31563)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_419.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[4]), .C(n31567), 
         .D(n31569), .Z(n29372)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21904_2_lut_rep_355_3_lut_4_lut (.A(state[1]), .B(state[4]), .C(uart_rx_c), 
         .D(n31569), .Z(n31499)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i21904_2_lut_rep_355_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_72 (.A(state[1]), .B(state[4]), .C(n31569), 
         .D(state[0]), .Z(n24509)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_3_lut_4_lut_adj_72.init = 16'hfffe;
    PFUMX i40 (.BLUT(n25), .ALUT(n27_adj_34), .C0(state[0]), .Z(n28399));
    LUT4 i14721_2_lut_rep_423 (.A(state[0]), .B(state[5]), .Z(n31567)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14721_2_lut_rep_423.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(state[0]), .B(state[5]), .C(state[4]), .Z(n13560)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_rep_424 (.A(state[1]), .B(bclk), .Z(n31568)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i1_2_lut_rep_424.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_adj_73 (.A(state[1]), .B(bclk), .C(state[3]), 
         .Z(n29384)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i1_2_lut_3_lut_adj_73.init = 16'hbfbf;
    LUT4 i2_2_lut_rep_425 (.A(state[3]), .B(state[2]), .Z(n31569)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_2_lut_rep_425.init = 16'heeee;
    LUT4 i1_2_lut_rep_376_3_lut_4_lut (.A(state[3]), .B(state[2]), .C(state[4]), 
         .D(state[1]), .Z(n31520)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_376_3_lut_4_lut.init = 16'hfffe;
    LUT4 state_1__bdd_2_lut (.A(state[1]), .B(bclk), .Z(n30709)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam state_1__bdd_2_lut.init = 16'h9999;
    PFUMX i36 (.BLUT(n21), .ALUT(n23), .C0(state[5]), .Z(n28051));
    PFUMX i9866 (.BLUT(n29203), .ALUT(n16637), .C0(state[0]), .Z(n16638));
    LUT4 state_1__bdd_4_lut (.A(state[1]), .B(n31519), .C(n31520), .D(uart_rx_c), 
         .Z(n30710)) /* synthesis lut_function=(A (B+!(C))+!A !(C+(D))) */ ;
    defparam state_1__bdd_4_lut.init = 16'h8a8f;
    LUT4 i41_4_lut_3_lut (.A(bclk), .B(state[1]), .C(state[2]), .Z(n27_adj_34)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i41_4_lut_3_lut.init = 16'hb4b4;
    LUT4 i1_4_lut_adj_74 (.A(rdata[0]), .B(rx_data[0]), .C(n13569), .D(n19_adj_32), 
         .Z(n9401)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_74.init = 16'heca0;
    FD1P3AX rdata_i0_i1 (.D(n9415), .SP(n31501), .CK(debug_c_c), .Q(rdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i1.GSR = "ENABLED";
    FD1P3AX rdata_i0_i2 (.D(n9417), .SP(n31501), .CK(debug_c_c), .Q(rdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i2.GSR = "ENABLED";
    FD1P3AX rdata_i0_i3 (.D(n9419), .SP(n31501), .CK(debug_c_c), .Q(rdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i3.GSR = "ENABLED";
    FD1P3AX rdata_i0_i4 (.D(n9421), .SP(n31501), .CK(debug_c_c), .Q(rdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i4.GSR = "ENABLED";
    FD1P3AX rdata_i0_i5 (.D(n9423), .SP(n31501), .CK(debug_c_c), .Q(rdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i5.GSR = "ENABLED";
    FD1P3AX rdata_i0_i6 (.D(n9425), .SP(n31501), .CK(debug_c_c), .Q(rdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i6.GSR = "ENABLED";
    FD1P3AX rdata_i0_i7 (.D(n9427), .SP(n31501), .CK(debug_c_c), .Q(rdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i7.GSR = "ENABLED";
    FD1P3AX data_i0_i1 (.D(n9429), .SP(n31501), .CK(debug_c_c), .Q(rx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i1.GSR = "ENABLED";
    FD1P3AX data_i0_i2 (.D(n9431), .SP(n31501), .CK(debug_c_c), .Q(rx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i2.GSR = "ENABLED";
    FD1P3AX data_i0_i3 (.D(n9433), .SP(n31501), .CK(debug_c_c), .Q(rx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i3.GSR = "ENABLED";
    FD1P3AX data_i0_i4 (.D(n9435), .SP(n31501), .CK(debug_c_c), .Q(rx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i4.GSR = "ENABLED";
    FD1P3AX data_i0_i5 (.D(n9437), .SP(n31501), .CK(debug_c_c), .Q(rx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i5.GSR = "ENABLED";
    FD1P3AX data_i0_i6 (.D(n9439), .SP(n31501), .CK(debug_c_c), .Q(rx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i6.GSR = "ENABLED";
    FD1P3AX data_i0_i7 (.D(n9441), .SP(n31501), .CK(debug_c_c), .Q(rx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i7.GSR = "ENABLED";
    FD1S3IX state__i1 (.D(n31404), .CK(debug_c_c), .CD(n31473), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i1.GSR = "ENABLED";
    FD1S3IX state__i2 (.D(n28399), .CK(debug_c_c), .CD(n31473), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i2.GSR = "ENABLED";
    FD1S3IX state__i3 (.D(n28297), .CK(debug_c_c), .CD(n31473), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i3.GSR = "ENABLED";
    FD1S3IX state__i4 (.D(n16638), .CK(debug_c_c), .CD(n31473), .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i4.GSR = "ENABLED";
    FD1S3IX state__i5 (.D(n28051), .CK(debug_c_c), .CD(n31473), .Q(state[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i5.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_75 (.A(state[5]), .B(n31499), .C(state[2]), .D(n31498), 
         .Z(n25)) /* synthesis lut_function=(!(A+!((C (D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_75.init = 16'h5111;
    LUT4 i15065_2_lut_rep_459 (.A(bclk), .B(state[1]), .Z(n31603)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15065_2_lut_rep_459.init = 16'h8888;
    LUT4 i15469_2_lut_3_lut (.A(bclk), .B(state[1]), .C(state[3]), .Z(n22201)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15469_2_lut_3_lut.init = 16'h8080;
    LUT4 i2_4_lut (.A(bclk), .B(n4), .C(state[0]), .D(n31519), .Z(n21)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i2_4_lut.init = 16'h4840;
    LUT4 i1_2_lut_adj_76 (.A(state[4]), .B(n10239), .Z(n4)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_76.init = 16'h8888;
    LUT4 i38_4_lut (.A(n31499), .B(n10239), .C(state[0]), .D(n4_adj_35), 
         .Z(n23)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i38_4_lut.init = 16'hf535;
    LUT4 i1_2_lut_adj_77 (.A(state[4]), .B(bclk), .Z(n4_adj_35)) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_77.init = 16'hdddd;
    LUT4 i22427_4_lut (.A(baud_reset), .B(n29372), .C(uart_rx_c), .D(n24509), 
         .Z(n19)) /* synthesis lut_function=(A (B+(C))+!A !((D)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i22427_4_lut.init = 16'ha8ec;
    LUT4 i3448_4_lut (.A(state[3]), .B(state[2]), .C(state[1]), .D(state[0]), 
         .Z(n10239)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3448_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_78 (.A(n78[0]), .B(rdata[0]), .C(n13560), .D(n13), 
         .Z(n9399)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_78.init = 16'heca0;
    LUT4 i4454_4_lut (.A(uart_rx_c), .B(rdata[0]), .C(n31569), .D(n31568), 
         .Z(n78[0])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4454_4_lut.init = 16'hccca;
    LUT4 i2_3_lut (.A(state[0]), .B(state[5]), .C(state[4]), .Z(n13)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_3_lut.init = 16'hefef;
    LUT4 rx_data_1__bdd_4_lut (.A(rx_data[1]), .B(rx_data[3]), .C(rx_data[4]), 
         .D(rx_data[2]), .Z(n30735)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C (D)))+!A (B+(C+(D)))) */ ;
    defparam rx_data_1__bdd_4_lut.init = 16'hdf7e;
    LUT4 i1_4_lut_adj_79 (.A(n1502), .B(debug_c_7), .C(n1504), .D(n51), 
         .Z(n13465)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_79.init = 16'heeea;
    LUT4 i47_4_lut (.A(n31454), .B(n1506), .C(n47), .D(n57), .Z(n51)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i47_4_lut.init = 16'h4f45;
    LUT4 i1_2_lut_adj_80 (.A(escape), .B(n1503), .Z(n47)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_80.init = 16'hbbbb;
    LUT4 i1_3_lut (.A(debug_c_7), .B(n1504), .C(n1503), .Z(n12482)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;
    defparam i1_3_lut.init = 16'h5454;
    LUT4 i1_2_lut_adj_81 (.A(rx_data[4]), .B(rx_data[3]), .Z(n29393)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_81.init = 16'heeee;
    \ClockDividerP(factor=12)_U0  baud_gen (.GND_net(GND_net), .baud_reset(baud_reset), 
            .bclk(bclk), .debug_c_c(debug_c_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(25[28] 27[56])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12)_U0 
//

module \ClockDividerP(factor=12)_U0  (GND_net, baud_reset, bclk, debug_c_c) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input baud_reset;
    output bclk;
    input debug_c_c;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26987;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n134;
    
    wire n26986, n26985, n26984, n26983, n26982, n26981, n26980, 
        n26979, n26978, n26977, n26976, n26975, n26974, n26973, 
        n26972, n57, n55, n56, n2963, n54, n46, n29624, n50, 
        n38, n52, n42, n48, n34, n8437, n27099, n27098, n27097, 
        n27096, n27095, n27094, n27093, n27092, n27091, n27090, 
        n27089, n27088, n27087, n27086, n27085, n27084;
    
    CCU2D count_2678_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26987), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_33.INIT1 = 16'h0000;
    defparam count_2678_add_4_33.INJECT1_0 = "NO";
    defparam count_2678_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26986), .COUT(n26987), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_31.INJECT1_0 = "NO";
    defparam count_2678_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26985), .COUT(n26986), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_29.INJECT1_0 = "NO";
    defparam count_2678_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26984), .COUT(n26985), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_27.INJECT1_0 = "NO";
    defparam count_2678_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26983), .COUT(n26984), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_25.INJECT1_0 = "NO";
    defparam count_2678_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26982), .COUT(n26983), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_23.INJECT1_0 = "NO";
    defparam count_2678_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26981), .COUT(n26982), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_21.INJECT1_0 = "NO";
    defparam count_2678_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26980), .COUT(n26981), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_19.INJECT1_0 = "NO";
    defparam count_2678_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26979), .COUT(n26980), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_17.INJECT1_0 = "NO";
    defparam count_2678_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26978), .COUT(n26979), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_15.INJECT1_0 = "NO";
    defparam count_2678_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26977), .COUT(n26978), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_13.INJECT1_0 = "NO";
    defparam count_2678_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26976), .COUT(n26977), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_11.INJECT1_0 = "NO";
    defparam count_2678_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26975), .COUT(n26976), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_9.INJECT1_0 = "NO";
    defparam count_2678_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26974), .COUT(n26975), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_7.INJECT1_0 = "NO";
    defparam count_2678_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26973), .COUT(n26974), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_5.INJECT1_0 = "NO";
    defparam count_2678_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26972), .COUT(n26973), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2678_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2678_add_4_3.INJECT1_0 = "NO";
    defparam count_2678_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2678_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26972), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678_add_4_1.INIT0 = 16'hF000;
    defparam count_2678_add_4_1.INIT1 = 16'h0555;
    defparam count_2678_add_4_1.INJECT1_0 = "NO";
    defparam count_2678_add_4_1.INJECT1_1 = "NO";
    LUT4 i1113_4_lut (.A(n57), .B(baud_reset), .C(n55), .D(n56), .Z(n2963)) /* synthesis lut_function=(A (B)+!A (B+!(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(23[5] 33[8])
    defparam i1113_4_lut.init = 16'hcccd;
    LUT4 i27_4_lut (.A(count[31]), .B(n54), .C(n46), .D(n29624), .Z(n57)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i27_4_lut.init = 16'hfeff;
    LUT4 i25_4_lut (.A(count[24]), .B(n50), .C(n38), .D(count[4]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(count[5]), .B(n52), .C(n42), .D(count[6]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(count[16]), .B(n48), .C(n34), .D(count[11]), 
         .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(count[28]), .B(count[2]), .C(count[18]), .D(count[8]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i22065_3_lut (.A(count[3]), .B(count[0]), .C(count[1]), .Z(n29624)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i22065_3_lut.init = 16'h8080;
    LUT4 i18_4_lut (.A(count[26]), .B(count[12]), .C(count[9]), .D(count[17]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(count[21]), .B(count[25]), .Z(n34)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i4_2_lut.init = 16'heeee;
    FD1S3IX clk_o_14 (.D(n8437), .CK(debug_c_c), .CD(baud_reset), .Q(bclk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    LUT4 i20_4_lut (.A(count[7]), .B(count[19]), .C(count[14]), .D(count[22]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(count[27]), .B(count[30]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i22_4_lut (.A(count[15]), .B(count[29]), .C(count[23]), .D(count[13]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i12_2_lut (.A(count[10]), .B(count[20]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i12_2_lut.init = 16'heeee;
    FD1S3IX count_2678__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2963), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i0.GSR = "ENABLED";
    CCU2D sub_2084_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27099), .S0(n8437));
    defparam sub_2084_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2084_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2084_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2084_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27098), .COUT(n27099));
    defparam sub_2084_add_2_32.INIT0 = 16'h5555;
    defparam sub_2084_add_2_32.INIT1 = 16'h5555;
    defparam sub_2084_add_2_32.INJECT1_0 = "NO";
    defparam sub_2084_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27097), .COUT(n27098));
    defparam sub_2084_add_2_30.INIT0 = 16'h5555;
    defparam sub_2084_add_2_30.INIT1 = 16'h5555;
    defparam sub_2084_add_2_30.INJECT1_0 = "NO";
    defparam sub_2084_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27096), .COUT(n27097));
    defparam sub_2084_add_2_28.INIT0 = 16'h5555;
    defparam sub_2084_add_2_28.INIT1 = 16'h5555;
    defparam sub_2084_add_2_28.INJECT1_0 = "NO";
    defparam sub_2084_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27095), .COUT(n27096));
    defparam sub_2084_add_2_26.INIT0 = 16'h5555;
    defparam sub_2084_add_2_26.INIT1 = 16'h5555;
    defparam sub_2084_add_2_26.INJECT1_0 = "NO";
    defparam sub_2084_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27094), .COUT(n27095));
    defparam sub_2084_add_2_24.INIT0 = 16'h5555;
    defparam sub_2084_add_2_24.INIT1 = 16'h5555;
    defparam sub_2084_add_2_24.INJECT1_0 = "NO";
    defparam sub_2084_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27093), .COUT(n27094));
    defparam sub_2084_add_2_22.INIT0 = 16'h5555;
    defparam sub_2084_add_2_22.INIT1 = 16'h5555;
    defparam sub_2084_add_2_22.INJECT1_0 = "NO";
    defparam sub_2084_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27092), .COUT(n27093));
    defparam sub_2084_add_2_20.INIT0 = 16'h5555;
    defparam sub_2084_add_2_20.INIT1 = 16'h5555;
    defparam sub_2084_add_2_20.INJECT1_0 = "NO";
    defparam sub_2084_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27091), .COUT(n27092));
    defparam sub_2084_add_2_18.INIT0 = 16'h5555;
    defparam sub_2084_add_2_18.INIT1 = 16'h5555;
    defparam sub_2084_add_2_18.INJECT1_0 = "NO";
    defparam sub_2084_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27090), .COUT(n27091));
    defparam sub_2084_add_2_16.INIT0 = 16'h5555;
    defparam sub_2084_add_2_16.INIT1 = 16'h5555;
    defparam sub_2084_add_2_16.INJECT1_0 = "NO";
    defparam sub_2084_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27089), .COUT(n27090));
    defparam sub_2084_add_2_14.INIT0 = 16'h5555;
    defparam sub_2084_add_2_14.INIT1 = 16'h5555;
    defparam sub_2084_add_2_14.INJECT1_0 = "NO";
    defparam sub_2084_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27088), .COUT(n27089));
    defparam sub_2084_add_2_12.INIT0 = 16'h5555;
    defparam sub_2084_add_2_12.INIT1 = 16'h5555;
    defparam sub_2084_add_2_12.INJECT1_0 = "NO";
    defparam sub_2084_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27087), .COUT(n27088));
    defparam sub_2084_add_2_10.INIT0 = 16'h5555;
    defparam sub_2084_add_2_10.INIT1 = 16'h5555;
    defparam sub_2084_add_2_10.INJECT1_0 = "NO";
    defparam sub_2084_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27086), .COUT(n27087));
    defparam sub_2084_add_2_8.INIT0 = 16'h5555;
    defparam sub_2084_add_2_8.INIT1 = 16'h5555;
    defparam sub_2084_add_2_8.INJECT1_0 = "NO";
    defparam sub_2084_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27085), .COUT(n27086));
    defparam sub_2084_add_2_6.INIT0 = 16'h5555;
    defparam sub_2084_add_2_6.INIT1 = 16'h5555;
    defparam sub_2084_add_2_6.INJECT1_0 = "NO";
    defparam sub_2084_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27084), .COUT(n27085));
    defparam sub_2084_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2084_add_2_4.INIT1 = 16'h5555;
    defparam sub_2084_add_2_4.INJECT1_0 = "NO";
    defparam sub_2084_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_2084_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27084));
    defparam sub_2084_add_2_2.INIT0 = 16'h0000;
    defparam sub_2084_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2084_add_2_2.INJECT1_0 = "NO";
    defparam sub_2084_add_2_2.INJECT1_1 = "NO";
    FD1S3IX count_2678__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2963), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i1.GSR = "ENABLED";
    FD1S3IX count_2678__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2963), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i2.GSR = "ENABLED";
    FD1S3IX count_2678__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2963), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i3.GSR = "ENABLED";
    FD1S3IX count_2678__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2963), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i4.GSR = "ENABLED";
    FD1S3IX count_2678__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2963), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i5.GSR = "ENABLED";
    FD1S3IX count_2678__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2963), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i6.GSR = "ENABLED";
    FD1S3IX count_2678__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2963), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i7.GSR = "ENABLED";
    FD1S3IX count_2678__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2963), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i8.GSR = "ENABLED";
    FD1S3IX count_2678__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2963), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i9.GSR = "ENABLED";
    FD1S3IX count_2678__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i10.GSR = "ENABLED";
    FD1S3IX count_2678__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i11.GSR = "ENABLED";
    FD1S3IX count_2678__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i12.GSR = "ENABLED";
    FD1S3IX count_2678__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i13.GSR = "ENABLED";
    FD1S3IX count_2678__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i14.GSR = "ENABLED";
    FD1S3IX count_2678__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i15.GSR = "ENABLED";
    FD1S3IX count_2678__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i16.GSR = "ENABLED";
    FD1S3IX count_2678__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i17.GSR = "ENABLED";
    FD1S3IX count_2678__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i18.GSR = "ENABLED";
    FD1S3IX count_2678__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i19.GSR = "ENABLED";
    FD1S3IX count_2678__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i20.GSR = "ENABLED";
    FD1S3IX count_2678__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i21.GSR = "ENABLED";
    FD1S3IX count_2678__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i22.GSR = "ENABLED";
    FD1S3IX count_2678__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i23.GSR = "ENABLED";
    FD1S3IX count_2678__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i24.GSR = "ENABLED";
    FD1S3IX count_2678__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i25.GSR = "ENABLED";
    FD1S3IX count_2678__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i26.GSR = "ENABLED";
    FD1S3IX count_2678__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i27.GSR = "ENABLED";
    FD1S3IX count_2678__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i28.GSR = "ENABLED";
    FD1S3IX count_2678__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i29.GSR = "ENABLED";
    FD1S3IX count_2678__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i30.GSR = "ENABLED";
    FD1S3IX count_2678__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2963), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2678__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module GlobalControlPeripheral
//

module GlobalControlPeripheral (\register[2] , GND_net, force_pause, debug_c_c, 
            n31512, \databus[1] , n9484, read_size, n14454, n31450, 
            prev_clk_1Hz, clk_1Hz, \register[0][2] , \select[1] , read_value, 
            n29069, rw, n46, n29293, n31478, n29294, n29295, n30306, 
            n30304, \reset_count[14] , n22484, xbee_pause_c, \register_addr[1] , 
            \register_addr[0] , n29170, n9538, n6003, n29066, n29056, 
            n29053, n16765, n27428, n29065, n16764, n29063, n29050, 
            n29052, n29054, n29067, n29057, n29068, n29071, n29072, 
            n29070, n6006, n29058, n29059, n29064, n29060, n29062, 
            n29055, n29051, n29049, n29061, n29048, n29789, n2876) /* synthesis syn_module_defined=1 */ ;
    output [31:0]\register[2] ;
    input GND_net;
    output force_pause;
    input debug_c_c;
    input n31512;
    input \databus[1] ;
    input n9484;
    output [2:0]read_size;
    output n14454;
    input n31450;
    output prev_clk_1Hz;
    output clk_1Hz;
    output \register[0][2] ;
    input \select[1] ;
    output [31:0]read_value;
    input n29069;
    input rw;
    output n46;
    input n29293;
    input n31478;
    input n29294;
    input n29295;
    input n30306;
    input n30304;
    input \reset_count[14] ;
    input n22484;
    input xbee_pause_c;
    input \register_addr[1] ;
    input \register_addr[0] ;
    output n29170;
    input n9538;
    input n6003;
    input n29066;
    input n29056;
    input n29053;
    input n16765;
    input n27428;
    input n29065;
    input n16764;
    input n29063;
    input n29050;
    input n29052;
    input n29054;
    input n29067;
    input n29057;
    input n29068;
    input n29071;
    input n29072;
    input n29070;
    input n6006;
    input n29058;
    input n29059;
    input n29064;
    input n29060;
    input n29062;
    input n29055;
    input n29051;
    input n29049;
    input n29061;
    input n29048;
    output n29789;
    input n2876;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26725;
    wire [31:0]n100;
    
    wire n26726, n26724, n26723, n26722, n27237, n26721, n179, 
        prev_select, n26720, n26719, n26718, n26717, n26716, n31592, 
        n26731, n26730, n26729, n26728, n26727;
    
    CCU2D add_135_21 (.A0(\register[2] [19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26725), .COUT(n26726), .S0(n100[19]), 
          .S1(n100[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_21.INIT0 = 16'h5aaa;
    defparam add_135_21.INIT1 = 16'h5aaa;
    defparam add_135_21.INJECT1_0 = "NO";
    defparam add_135_21.INJECT1_1 = "NO";
    CCU2D add_135_19 (.A0(\register[2] [17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26724), .COUT(n26725), .S0(n100[17]), 
          .S1(n100[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_19.INIT0 = 16'h5aaa;
    defparam add_135_19.INIT1 = 16'h5aaa;
    defparam add_135_19.INJECT1_0 = "NO";
    defparam add_135_19.INJECT1_1 = "NO";
    CCU2D add_135_17 (.A0(\register[2] [15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26723), .COUT(n26724), .S0(n100[15]), 
          .S1(n100[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_17.INIT0 = 16'h5aaa;
    defparam add_135_17.INIT1 = 16'h5aaa;
    defparam add_135_17.INJECT1_0 = "NO";
    defparam add_135_17.INJECT1_1 = "NO";
    CCU2D add_135_15 (.A0(\register[2] [13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26722), .COUT(n26723), .S0(n100[13]), 
          .S1(n100[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_15.INIT0 = 16'h5aaa;
    defparam add_135_15.INIT1 = 16'h5aaa;
    defparam add_135_15.INJECT1_0 = "NO";
    defparam add_135_15.INJECT1_1 = "NO";
    FD1P3IX force_pause_152 (.D(\databus[1] ), .SP(n27237), .CD(n31512), 
            .CK(debug_c_c), .Q(force_pause));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam force_pause_152.GSR = "ENABLED";
    CCU2D add_135_13 (.A0(\register[2] [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26721), .COUT(n26722), .S0(n100[11]), 
          .S1(n100[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_13.INIT0 = 16'h5aaa;
    defparam add_135_13.INIT1 = 16'h5aaa;
    defparam add_135_13.INJECT1_0 = "NO";
    defparam add_135_13.INJECT1_1 = "NO";
    FD1P3IX uptime_count__i31 (.D(n100[31]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i31.GSR = "ENABLED";
    FD1P3IX uptime_count__i30 (.D(n100[30]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i30.GSR = "ENABLED";
    FD1P3IX uptime_count__i29 (.D(n100[29]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i29.GSR = "ENABLED";
    FD1P3IX uptime_count__i28 (.D(n100[28]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i28.GSR = "ENABLED";
    FD1P3IX uptime_count__i27 (.D(n100[27]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i27.GSR = "ENABLED";
    FD1P3IX uptime_count__i26 (.D(n100[26]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i26.GSR = "ENABLED";
    FD1P3IX uptime_count__i25 (.D(n100[25]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i25.GSR = "ENABLED";
    FD1P3IX uptime_count__i24 (.D(n100[24]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i24.GSR = "ENABLED";
    FD1P3IX uptime_count__i23 (.D(n100[23]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i23.GSR = "ENABLED";
    FD1P3IX uptime_count__i22 (.D(n100[22]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i22.GSR = "ENABLED";
    FD1P3IX uptime_count__i21 (.D(n100[21]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i21.GSR = "ENABLED";
    FD1P3IX uptime_count__i20 (.D(n100[20]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i20.GSR = "ENABLED";
    FD1P3IX uptime_count__i19 (.D(n100[19]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i19.GSR = "ENABLED";
    FD1P3IX uptime_count__i18 (.D(n100[18]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i18.GSR = "ENABLED";
    FD1P3IX uptime_count__i17 (.D(n100[17]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i17.GSR = "ENABLED";
    FD1P3IX uptime_count__i16 (.D(n100[16]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i16.GSR = "ENABLED";
    FD1P3IX uptime_count__i15 (.D(n100[15]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i15.GSR = "ENABLED";
    FD1P3IX uptime_count__i14 (.D(n100[14]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i14.GSR = "ENABLED";
    FD1P3IX uptime_count__i13 (.D(n100[13]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i13.GSR = "ENABLED";
    FD1P3IX uptime_count__i12 (.D(n100[12]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i12.GSR = "ENABLED";
    FD1P3IX uptime_count__i11 (.D(n100[11]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i11.GSR = "ENABLED";
    FD1P3IX uptime_count__i10 (.D(n100[10]), .SP(n9484), .CD(n31512), 
            .CK(debug_c_c), .Q(\register[2] [10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i10.GSR = "ENABLED";
    FD1P3IX uptime_count__i9 (.D(n100[9]), .SP(n9484), .CD(n31512), .CK(debug_c_c), 
            .Q(\register[2] [9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i9.GSR = "ENABLED";
    FD1P3IX uptime_count__i8 (.D(n100[8]), .SP(n9484), .CD(n31512), .CK(debug_c_c), 
            .Q(\register[2] [8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i8.GSR = "ENABLED";
    FD1P3IX uptime_count__i7 (.D(n100[7]), .SP(n9484), .CD(n31512), .CK(debug_c_c), 
            .Q(\register[2] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i7.GSR = "ENABLED";
    FD1P3IX uptime_count__i6 (.D(n100[6]), .SP(n9484), .CD(n31512), .CK(debug_c_c), 
            .Q(\register[2] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i6.GSR = "ENABLED";
    FD1P3IX uptime_count__i5 (.D(n100[5]), .SP(n9484), .CD(n31512), .CK(debug_c_c), 
            .Q(\register[2] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i5.GSR = "ENABLED";
    FD1P3IX uptime_count__i4 (.D(n100[4]), .SP(n9484), .CD(n31512), .CK(debug_c_c), 
            .Q(\register[2] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i4.GSR = "ENABLED";
    FD1P3IX uptime_count__i3 (.D(n100[3]), .SP(n9484), .CD(n31512), .CK(debug_c_c), 
            .Q(\register[2] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i3.GSR = "ENABLED";
    FD1P3IX uptime_count__i2 (.D(n100[2]), .SP(n9484), .CD(n31512), .CK(debug_c_c), 
            .Q(\register[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i2.GSR = "ENABLED";
    FD1P3IX uptime_count__i1 (.D(n100[1]), .SP(n9484), .CD(n31512), .CK(debug_c_c), 
            .Q(\register[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i1.GSR = "ENABLED";
    FD1P3IX uptime_count__i0 (.D(n100[0]), .SP(n9484), .CD(n31512), .CK(debug_c_c), 
            .Q(\register[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i0.GSR = "ENABLED";
    FD1P3AX read_size_i0_i0 (.D(n31450), .SP(n14454), .CK(debug_c_c), 
            .Q(read_size[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_size_i0_i0.GSR = "ENABLED";
    FD1S3AX prev_clk_1Hz_150 (.D(clk_1Hz), .CK(debug_c_c), .Q(prev_clk_1Hz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam prev_clk_1Hz_150.GSR = "ENABLED";
    FD1S3AX xbee_pause_latched_151 (.D(n179), .CK(debug_c_c), .Q(\register[0][2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam xbee_pause_latched_151.GSR = "ENABLED";
    FD1S3AX prev_select_149 (.D(\select[1] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam prev_select_149.GSR = "ENABLED";
    CCU2D add_135_11 (.A0(\register[2] [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26720), .COUT(n26721), .S0(n100[9]), .S1(n100[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_11.INIT0 = 16'h5aaa;
    defparam add_135_11.INIT1 = 16'h5aaa;
    defparam add_135_11.INJECT1_0 = "NO";
    defparam add_135_11.INJECT1_1 = "NO";
    CCU2D add_135_9 (.A0(\register[2] [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26719), .COUT(n26720), .S0(n100[7]), .S1(n100[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_9.INIT0 = 16'h5aaa;
    defparam add_135_9.INIT1 = 16'h5aaa;
    defparam add_135_9.INJECT1_0 = "NO";
    defparam add_135_9.INJECT1_1 = "NO";
    CCU2D add_135_7 (.A0(\register[2] [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26718), .COUT(n26719), .S0(n100[5]), .S1(n100[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_7.INIT0 = 16'h5aaa;
    defparam add_135_7.INIT1 = 16'h5aaa;
    defparam add_135_7.INJECT1_0 = "NO";
    defparam add_135_7.INJECT1_1 = "NO";
    CCU2D add_135_5 (.A0(\register[2] [3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26717), .COUT(n26718), .S0(n100[3]), .S1(n100[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_5.INIT0 = 16'h5aaa;
    defparam add_135_5.INIT1 = 16'h5aaa;
    defparam add_135_5.INJECT1_0 = "NO";
    defparam add_135_5.INJECT1_1 = "NO";
    CCU2D add_135_3 (.A0(\register[2] [1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26716), .COUT(n26717), .S0(n100[1]), .S1(n100[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_3.INIT0 = 16'h5aaa;
    defparam add_135_3.INIT1 = 16'h5aaa;
    defparam add_135_3.INJECT1_0 = "NO";
    defparam add_135_3.INJECT1_1 = "NO";
    CCU2D add_135_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\register[2] [0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26716), .S1(n100[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_1.INIT0 = 16'hF000;
    defparam add_135_1.INIT1 = 16'h5555;
    defparam add_135_1.INJECT1_0 = "NO";
    defparam add_135_1.INJECT1_1 = "NO";
    FD1P3AX read_value__i28 (.D(n29069), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i28.GSR = "ENABLED";
    LUT4 i14_2_lut (.A(\select[1] ), .B(rw), .Z(n46)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(36[19:32])
    defparam i14_2_lut.init = 16'h8888;
    FD1P3AX read_value__i29 (.D(n29293), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i29.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(n31512), .B(rw), .C(n31592), .D(n31478), .Z(n27237)) /* synthesis lut_function=(!(A (B+(D))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam i2_4_lut.init = 16'h0032;
    FD1P3AX read_value__i30 (.D(n29294), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n29295), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX read_value__i2 (.D(n30306), .SP(n14454), .CK(debug_c_c), .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3AX read_value__i1 (.D(n30304), .SP(n14454), .CK(debug_c_c), .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i118_2_lut_rep_448 (.A(prev_select), .B(\select[1] ), .Z(n31592)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(60[9:30])
    defparam i118_2_lut_rep_448.init = 16'h4444;
    LUT4 i965_2_lut_2_lut_3_lut_4_lut (.A(prev_select), .B(\select[1] ), 
         .C(\reset_count[14] ), .D(n22484), .Z(n14454)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(60[9:30])
    defparam i965_2_lut_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i115_1_lut (.A(xbee_pause_c), .Z(n179)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(52[26:39])
    defparam i115_1_lut.init = 16'h5555;
    LUT4 i1_2_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), .Z(n29170)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut.init = 16'h2222;
    FD1P3IX read_value__i3 (.D(n6003), .SP(n14454), .CD(n9538), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3AX read_value__i4 (.D(n29066), .SP(n14454), .CK(debug_c_c), .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3AX read_value__i5 (.D(n29056), .SP(n14454), .CK(debug_c_c), .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3AX read_value__i6 (.D(n29053), .SP(n14454), .CK(debug_c_c), .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_size_i0_i1 (.D(n27428), .SP(n14454), .CD(n16765), .CK(debug_c_c), 
            .Q(read_size[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_size_i0_i1.GSR = "ENABLED";
    FD1P3AX read_value__i7 (.D(n29065), .SP(n14454), .CK(debug_c_c), .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_size_i0_i2 (.D(n31478), .SP(n14454), .CD(n16764), .CK(debug_c_c), 
            .Q(read_size[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_size_i0_i2.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29063), .SP(n14454), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29050), .SP(n14454), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29052), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29054), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29067), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29057), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29068), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29071), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29072), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29070), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n6006), .SP(n14454), .CD(n9538), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29058), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n29059), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29064), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29060), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29062), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29055), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29051), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i24.GSR = "ENABLED";
    CCU2D add_135_33 (.A0(\register[2] [31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26731), .S0(n100[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_33.INIT0 = 16'h5aaa;
    defparam add_135_33.INIT1 = 16'h0000;
    defparam add_135_33.INJECT1_0 = "NO";
    defparam add_135_33.INJECT1_1 = "NO";
    CCU2D add_135_31 (.A0(\register[2] [29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26730), .COUT(n26731), .S0(n100[29]), 
          .S1(n100[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_31.INIT0 = 16'h5aaa;
    defparam add_135_31.INIT1 = 16'h5aaa;
    defparam add_135_31.INJECT1_0 = "NO";
    defparam add_135_31.INJECT1_1 = "NO";
    FD1P3AX read_value__i25 (.D(n29049), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i25.GSR = "ENABLED";
    CCU2D add_135_29 (.A0(\register[2] [27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26729), .COUT(n26730), .S0(n100[27]), 
          .S1(n100[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_29.INIT0 = 16'h5aaa;
    defparam add_135_29.INIT1 = 16'h5aaa;
    defparam add_135_29.INJECT1_0 = "NO";
    defparam add_135_29.INJECT1_1 = "NO";
    CCU2D add_135_27 (.A0(\register[2] [25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26728), .COUT(n26729), .S0(n100[25]), 
          .S1(n100[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_27.INIT0 = 16'h5aaa;
    defparam add_135_27.INIT1 = 16'h5aaa;
    defparam add_135_27.INJECT1_0 = "NO";
    defparam add_135_27.INJECT1_1 = "NO";
    CCU2D add_135_25 (.A0(\register[2] [23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26727), .COUT(n26728), .S0(n100[23]), 
          .S1(n100[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_25.INIT0 = 16'h5aaa;
    defparam add_135_25.INIT1 = 16'h5aaa;
    defparam add_135_25.INJECT1_0 = "NO";
    defparam add_135_25.INJECT1_1 = "NO";
    FD1P3AX read_value__i26 (.D(n29061), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i26.GSR = "ENABLED";
    CCU2D add_135_23 (.A0(\register[2] [21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26726), .COUT(n26727), .S0(n100[21]), 
          .S1(n100[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_23.INIT0 = 16'h5aaa;
    defparam add_135_23.INIT1 = 16'h5aaa;
    defparam add_135_23.INJECT1_0 = "NO";
    defparam add_135_23.INJECT1_1 = "NO";
    FD1P3AX read_value__i27 (.D(n29048), .SP(n14454), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i27.GSR = "ENABLED";
    \ClockDividerP(factor=12000000)  uptime_div (.GND_net(GND_net), .clk_1Hz(clk_1Hz), 
            .debug_c_c(debug_c_c), .n31512(n31512), .n29789(n29789), .n2876(n2876)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(105[28] 107[53])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000000) 
//

module \ClockDividerP(factor=12000000)  (GND_net, clk_1Hz, debug_c_c, 
            n31512, n29789, n2876) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output clk_1Hz;
    input debug_c_c;
    input n31512;
    output n29789;
    input n2876;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27181, n7986, n27180;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n27179, n27178, n27177, n27176, n27175, n27174, n27173, 
        n27172, n27171, n27170, n26971;
    wire [31:0]n134;
    
    wire n26970, n26969, n26968, n26967, n26966, n26965, n26964, 
        n26963, n26962, n26961, n26960, n26959, n26958, n26957, 
        n27, n27374, n25, n26, n24, n19, n32, n28, n20, n29, 
        n26_adj_30, n26956;
    
    CCU2D add_19624_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27181), 
          .S0(n7986));
    defparam add_19624_cout.INIT0 = 16'h0000;
    defparam add_19624_cout.INIT1 = 16'h0000;
    defparam add_19624_cout.INJECT1_0 = "NO";
    defparam add_19624_cout.INJECT1_1 = "NO";
    CCU2D add_19624_24 (.A0(count[30]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[31]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27180), .COUT(n27181));
    defparam add_19624_24.INIT0 = 16'h5555;
    defparam add_19624_24.INIT1 = 16'h5555;
    defparam add_19624_24.INJECT1_0 = "NO";
    defparam add_19624_24.INJECT1_1 = "NO";
    CCU2D add_19624_22 (.A0(count[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[29]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27179), .COUT(n27180));
    defparam add_19624_22.INIT0 = 16'h5555;
    defparam add_19624_22.INIT1 = 16'h5555;
    defparam add_19624_22.INJECT1_0 = "NO";
    defparam add_19624_22.INJECT1_1 = "NO";
    CCU2D add_19624_20 (.A0(count[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27178), .COUT(n27179));
    defparam add_19624_20.INIT0 = 16'h5555;
    defparam add_19624_20.INIT1 = 16'h5555;
    defparam add_19624_20.INJECT1_0 = "NO";
    defparam add_19624_20.INJECT1_1 = "NO";
    CCU2D add_19624_18 (.A0(count[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27177), .COUT(n27178));
    defparam add_19624_18.INIT0 = 16'h5555;
    defparam add_19624_18.INIT1 = 16'h5555;
    defparam add_19624_18.INJECT1_0 = "NO";
    defparam add_19624_18.INJECT1_1 = "NO";
    CCU2D add_19624_16 (.A0(count[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27176), .COUT(n27177));
    defparam add_19624_16.INIT0 = 16'h5aaa;
    defparam add_19624_16.INIT1 = 16'h5555;
    defparam add_19624_16.INJECT1_0 = "NO";
    defparam add_19624_16.INJECT1_1 = "NO";
    CCU2D add_19624_14 (.A0(count[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27175), .COUT(n27176));
    defparam add_19624_14.INIT0 = 16'h5aaa;
    defparam add_19624_14.INIT1 = 16'h5555;
    defparam add_19624_14.INJECT1_0 = "NO";
    defparam add_19624_14.INJECT1_1 = "NO";
    CCU2D add_19624_12 (.A0(count[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27174), .COUT(n27175));
    defparam add_19624_12.INIT0 = 16'h5555;
    defparam add_19624_12.INIT1 = 16'h5aaa;
    defparam add_19624_12.INJECT1_0 = "NO";
    defparam add_19624_12.INJECT1_1 = "NO";
    CCU2D add_19624_10 (.A0(count[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27173), .COUT(n27174));
    defparam add_19624_10.INIT0 = 16'h5aaa;
    defparam add_19624_10.INIT1 = 16'h5aaa;
    defparam add_19624_10.INJECT1_0 = "NO";
    defparam add_19624_10.INJECT1_1 = "NO";
    CCU2D add_19624_8 (.A0(count[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27172), .COUT(n27173));
    defparam add_19624_8.INIT0 = 16'h5555;
    defparam add_19624_8.INIT1 = 16'h5aaa;
    defparam add_19624_8.INJECT1_0 = "NO";
    defparam add_19624_8.INJECT1_1 = "NO";
    CCU2D add_19624_6 (.A0(count[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27171), .COUT(n27172));
    defparam add_19624_6.INIT0 = 16'h5555;
    defparam add_19624_6.INIT1 = 16'h5555;
    defparam add_19624_6.INJECT1_0 = "NO";
    defparam add_19624_6.INJECT1_1 = "NO";
    CCU2D add_19624_4 (.A0(count[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27170), .COUT(n27171));
    defparam add_19624_4.INIT0 = 16'h5aaa;
    defparam add_19624_4.INIT1 = 16'h5aaa;
    defparam add_19624_4.INJECT1_0 = "NO";
    defparam add_19624_4.INJECT1_1 = "NO";
    CCU2D add_19624_2 (.A0(count[8]), .B0(count[7]), .C0(GND_net), .D0(GND_net), 
          .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27170));
    defparam add_19624_2.INIT0 = 16'h7000;
    defparam add_19624_2.INIT1 = 16'h5555;
    defparam add_19624_2.INJECT1_0 = "NO";
    defparam add_19624_2.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26971), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_33.INIT1 = 16'h0000;
    defparam count_2673_add_4_33.INJECT1_0 = "NO";
    defparam count_2673_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26970), .COUT(n26971), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_31.INJECT1_0 = "NO";
    defparam count_2673_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26969), .COUT(n26970), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_29.INJECT1_0 = "NO";
    defparam count_2673_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26968), .COUT(n26969), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_27.INJECT1_0 = "NO";
    defparam count_2673_add_4_27.INJECT1_1 = "NO";
    FD1S3IX clk_o_14 (.D(n7986), .CK(debug_c_c), .CD(n31512), .Q(clk_1Hz));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D count_2673_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26967), .COUT(n26968), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_25.INJECT1_0 = "NO";
    defparam count_2673_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26966), .COUT(n26967), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_23.INJECT1_0 = "NO";
    defparam count_2673_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26965), .COUT(n26966), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_21.INJECT1_0 = "NO";
    defparam count_2673_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26964), .COUT(n26965), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_19.INJECT1_0 = "NO";
    defparam count_2673_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26963), .COUT(n26964), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_17.INJECT1_0 = "NO";
    defparam count_2673_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26962), .COUT(n26963), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_15.INJECT1_0 = "NO";
    defparam count_2673_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26961), .COUT(n26962), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_13.INJECT1_0 = "NO";
    defparam count_2673_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26960), .COUT(n26961), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_11.INJECT1_0 = "NO";
    defparam count_2673_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26959), .COUT(n26960), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_9.INJECT1_0 = "NO";
    defparam count_2673_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26958), .COUT(n26959), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_7.INJECT1_0 = "NO";
    defparam count_2673_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2673_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26957), .COUT(n26958), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_5.INJECT1_0 = "NO";
    defparam count_2673_add_4_5.INJECT1_1 = "NO";
    LUT4 i22329_4_lut (.A(n27), .B(n27374), .C(n25), .D(n26), .Z(n29789)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i22329_4_lut.init = 16'h0004;
    LUT4 i12_4_lut (.A(count[19]), .B(n24), .C(count[8]), .D(count[14]), 
         .Z(n27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(n19), .B(n32), .C(n28), .D(n20), .Z(n27374)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16_4_lut.init = 16'h8000;
    LUT4 i10_4_lut (.A(count[30]), .B(count[22]), .C(count[13]), .D(count[25]), 
         .Z(n25)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i11_4_lut (.A(count[28]), .B(count[15]), .C(count[31]), .D(count[29]), 
         .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut (.A(count[26]), .B(count[24]), .C(count[10]), .D(count[27]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[18]), .B(count[1]), .Z(n19)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i15_4_lut (.A(n29), .B(count[9]), .C(n26_adj_30), .D(count[0]), 
         .Z(n32)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i15_4_lut.init = 16'h8000;
    LUT4 i11_4_lut_adj_55 (.A(count[3]), .B(count[12]), .C(count[5]), 
         .D(count[17]), .Z(n28)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i11_4_lut_adj_55.init = 16'h8000;
    LUT4 i3_2_lut (.A(count[2]), .B(count[11]), .Z(n20)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    CCU2D count_2673_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26956), .COUT(n26957), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2673_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2673_add_4_3.INJECT1_0 = "NO";
    defparam count_2673_add_4_3.INJECT1_1 = "NO";
    LUT4 i12_4_lut_adj_56 (.A(count[20]), .B(count[7]), .C(count[23]), 
         .D(count[21]), .Z(n29)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12_4_lut_adj_56.init = 16'h8000;
    CCU2D count_2673_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26956), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673_add_4_1.INIT0 = 16'hF000;
    defparam count_2673_add_4_1.INIT1 = 16'h0555;
    defparam count_2673_add_4_1.INJECT1_0 = "NO";
    defparam count_2673_add_4_1.INJECT1_1 = "NO";
    LUT4 i9_3_lut (.A(count[16]), .B(count[4]), .C(count[6]), .Z(n26_adj_30)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i9_3_lut.init = 16'h8080;
    FD1S3IX count_2673__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2876), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i0.GSR = "ENABLED";
    FD1S3IX count_2673__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2876), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i1.GSR = "ENABLED";
    FD1S3IX count_2673__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2876), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i2.GSR = "ENABLED";
    FD1S3IX count_2673__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2876), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i3.GSR = "ENABLED";
    FD1S3IX count_2673__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2876), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i4.GSR = "ENABLED";
    FD1S3IX count_2673__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2876), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i5.GSR = "ENABLED";
    FD1S3IX count_2673__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2876), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i6.GSR = "ENABLED";
    FD1S3IX count_2673__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2876), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i7.GSR = "ENABLED";
    FD1S3IX count_2673__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2876), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i8.GSR = "ENABLED";
    FD1S3IX count_2673__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2876), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i9.GSR = "ENABLED";
    FD1S3IX count_2673__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i10.GSR = "ENABLED";
    FD1S3IX count_2673__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i11.GSR = "ENABLED";
    FD1S3IX count_2673__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i12.GSR = "ENABLED";
    FD1S3IX count_2673__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i13.GSR = "ENABLED";
    FD1S3IX count_2673__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i14.GSR = "ENABLED";
    FD1S3IX count_2673__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i15.GSR = "ENABLED";
    FD1S3IX count_2673__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i16.GSR = "ENABLED";
    FD1S3IX count_2673__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i17.GSR = "ENABLED";
    FD1S3IX count_2673__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i18.GSR = "ENABLED";
    FD1S3IX count_2673__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i19.GSR = "ENABLED";
    FD1S3IX count_2673__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i20.GSR = "ENABLED";
    FD1S3IX count_2673__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i21.GSR = "ENABLED";
    FD1S3IX count_2673__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i22.GSR = "ENABLED";
    FD1S3IX count_2673__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i23.GSR = "ENABLED";
    FD1S3IX count_2673__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i24.GSR = "ENABLED";
    FD1S3IX count_2673__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i25.GSR = "ENABLED";
    FD1S3IX count_2673__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i26.GSR = "ENABLED";
    FD1S3IX count_2673__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i27.GSR = "ENABLED";
    FD1S3IX count_2673__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i28.GSR = "ENABLED";
    FD1S3IX count_2673__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i29.GSR = "ENABLED";
    FD1S3IX count_2673__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i30.GSR = "ENABLED";
    FD1S3IX count_2673__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2876), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2673__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module ClockDivider_U10
//

module ClockDivider_U10 (clk_255kHz, debug_c_c, n241, GND_net, n7917, 
            n31512, n7882, n29832, n14513, n29830, n14514, n2824, 
            n29840, n27541, n29847, n27536, n29818, n13957, n29530, 
            n14, n29944, n14500, n29784, n27564, n29811, n27547, 
            n29827, n27543, n29838, n27550) /* synthesis syn_module_defined=1 */ ;
    output clk_255kHz;
    input debug_c_c;
    input n241;
    input GND_net;
    output n7917;
    input n31512;
    output n7882;
    input n29832;
    output n14513;
    input n29830;
    output n14514;
    input n2824;
    input n29840;
    output n27541;
    input n29847;
    output n27536;
    input n29818;
    output n13957;
    input n29530;
    output n14;
    input n29944;
    output n14500;
    input n29784;
    output n27564;
    input n29811;
    output n27547;
    input n29827;
    output n27543;
    input n29838;
    output n27550;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26715, n26714;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    
    wire n26713, n26712, n26711, n26710, n26709, n26708, n26707, 
        n26706, n26705, n26704, n26703, n26702, n26701, n26700;
    wire [31:0]n134;
    
    wire n27130, n27129, n27128, n27127, n27126, n27125, n27124, 
        n27123, n27122, n27121, n27120, n27119, n27118, n27117, 
        n27116, n26907, n26906, n26905, n26904, n26903, n26902, 
        n26901, n26900, n26899, n26898, n26897, n26896, n26895, 
        n26894, n26893, n26892;
    
    FD1S3AX clk_o_22 (.D(n241), .CK(debug_c_c), .Q(clk_255kHz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=540, LSE_RLINE=543 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2059_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26715), .S0(n7917));
    defparam sub_2059_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2059_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2059_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2059_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26714), .COUT(n26715));
    defparam sub_2059_add_2_32.INIT0 = 16'h5555;
    defparam sub_2059_add_2_32.INIT1 = 16'h5555;
    defparam sub_2059_add_2_32.INJECT1_0 = "NO";
    defparam sub_2059_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26713), .COUT(n26714));
    defparam sub_2059_add_2_30.INIT0 = 16'h5555;
    defparam sub_2059_add_2_30.INIT1 = 16'h5555;
    defparam sub_2059_add_2_30.INJECT1_0 = "NO";
    defparam sub_2059_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26712), .COUT(n26713));
    defparam sub_2059_add_2_28.INIT0 = 16'h5555;
    defparam sub_2059_add_2_28.INIT1 = 16'h5555;
    defparam sub_2059_add_2_28.INJECT1_0 = "NO";
    defparam sub_2059_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26711), .COUT(n26712));
    defparam sub_2059_add_2_26.INIT0 = 16'h5555;
    defparam sub_2059_add_2_26.INIT1 = 16'h5555;
    defparam sub_2059_add_2_26.INJECT1_0 = "NO";
    defparam sub_2059_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26710), .COUT(n26711));
    defparam sub_2059_add_2_24.INIT0 = 16'h5555;
    defparam sub_2059_add_2_24.INIT1 = 16'h5555;
    defparam sub_2059_add_2_24.INJECT1_0 = "NO";
    defparam sub_2059_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26709), .COUT(n26710));
    defparam sub_2059_add_2_22.INIT0 = 16'h5555;
    defparam sub_2059_add_2_22.INIT1 = 16'h5555;
    defparam sub_2059_add_2_22.INJECT1_0 = "NO";
    defparam sub_2059_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26708), .COUT(n26709));
    defparam sub_2059_add_2_20.INIT0 = 16'h5555;
    defparam sub_2059_add_2_20.INIT1 = 16'h5555;
    defparam sub_2059_add_2_20.INJECT1_0 = "NO";
    defparam sub_2059_add_2_20.INJECT1_1 = "NO";
    LUT4 i22373_2_lut_4_lut (.A(n31512), .B(clk_255kHz), .C(n7882), .D(n29832), 
         .Z(n14513)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22373_2_lut_4_lut.init = 16'h1000;
    LUT4 i22371_2_lut_4_lut (.A(n31512), .B(clk_255kHz), .C(n7882), .D(n29830), 
         .Z(n14514)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22371_2_lut_4_lut.init = 16'h1000;
    CCU2D sub_2059_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26707), .COUT(n26708));
    defparam sub_2059_add_2_18.INIT0 = 16'h5555;
    defparam sub_2059_add_2_18.INIT1 = 16'h5555;
    defparam sub_2059_add_2_18.INJECT1_0 = "NO";
    defparam sub_2059_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26706), .COUT(n26707));
    defparam sub_2059_add_2_16.INIT0 = 16'h5555;
    defparam sub_2059_add_2_16.INIT1 = 16'h5555;
    defparam sub_2059_add_2_16.INJECT1_0 = "NO";
    defparam sub_2059_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26705), .COUT(n26706));
    defparam sub_2059_add_2_14.INIT0 = 16'h5555;
    defparam sub_2059_add_2_14.INIT1 = 16'h5555;
    defparam sub_2059_add_2_14.INJECT1_0 = "NO";
    defparam sub_2059_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26704), .COUT(n26705));
    defparam sub_2059_add_2_12.INIT0 = 16'h5555;
    defparam sub_2059_add_2_12.INIT1 = 16'h5555;
    defparam sub_2059_add_2_12.INJECT1_0 = "NO";
    defparam sub_2059_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26703), .COUT(n26704));
    defparam sub_2059_add_2_10.INIT0 = 16'h5555;
    defparam sub_2059_add_2_10.INIT1 = 16'h5555;
    defparam sub_2059_add_2_10.INJECT1_0 = "NO";
    defparam sub_2059_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26702), .COUT(n26703));
    defparam sub_2059_add_2_8.INIT0 = 16'h5555;
    defparam sub_2059_add_2_8.INIT1 = 16'h5555;
    defparam sub_2059_add_2_8.INJECT1_0 = "NO";
    defparam sub_2059_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26701), .COUT(n26702));
    defparam sub_2059_add_2_6.INIT0 = 16'h5555;
    defparam sub_2059_add_2_6.INIT1 = 16'h5aaa;
    defparam sub_2059_add_2_6.INJECT1_0 = "NO";
    defparam sub_2059_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26700), .COUT(n26701));
    defparam sub_2059_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2059_add_2_4.INIT1 = 16'h5aaa;
    defparam sub_2059_add_2_4.INJECT1_0 = "NO";
    defparam sub_2059_add_2_4.INJECT1_1 = "NO";
    FD1S3IX count_2671__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2824), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i0.GSR = "ENABLED";
    CCU2D sub_2059_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26700));
    defparam sub_2059_add_2_2.INIT0 = 16'h0000;
    defparam sub_2059_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2059_add_2_2.INJECT1_0 = "NO";
    defparam sub_2059_add_2_2.INJECT1_1 = "NO";
    LUT4 i22381_2_lut_4_lut (.A(n31512), .B(clk_255kHz), .C(n7882), .D(n29840), 
         .Z(n27541)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22381_2_lut_4_lut.init = 16'h1000;
    CCU2D add_19627_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27130), 
          .S1(n7882));
    defparam add_19627_32.INIT0 = 16'h5555;
    defparam add_19627_32.INIT1 = 16'h0000;
    defparam add_19627_32.INJECT1_0 = "NO";
    defparam add_19627_32.INJECT1_1 = "NO";
    CCU2D add_19627_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27129), .COUT(n27130));
    defparam add_19627_30.INIT0 = 16'h5555;
    defparam add_19627_30.INIT1 = 16'h5555;
    defparam add_19627_30.INJECT1_0 = "NO";
    defparam add_19627_30.INJECT1_1 = "NO";
    CCU2D add_19627_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27128), .COUT(n27129));
    defparam add_19627_28.INIT0 = 16'h5555;
    defparam add_19627_28.INIT1 = 16'h5555;
    defparam add_19627_28.INJECT1_0 = "NO";
    defparam add_19627_28.INJECT1_1 = "NO";
    CCU2D add_19627_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27127), .COUT(n27128));
    defparam add_19627_26.INIT0 = 16'h5555;
    defparam add_19627_26.INIT1 = 16'h5555;
    defparam add_19627_26.INJECT1_0 = "NO";
    defparam add_19627_26.INJECT1_1 = "NO";
    LUT4 i22388_2_lut_4_lut (.A(n31512), .B(clk_255kHz), .C(n7882), .D(n29847), 
         .Z(n27536)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22388_2_lut_4_lut.init = 16'h1000;
    CCU2D add_19627_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27126), .COUT(n27127));
    defparam add_19627_24.INIT0 = 16'h5555;
    defparam add_19627_24.INIT1 = 16'h5555;
    defparam add_19627_24.INJECT1_0 = "NO";
    defparam add_19627_24.INJECT1_1 = "NO";
    LUT4 i22359_2_lut_4_lut (.A(n31512), .B(clk_255kHz), .C(n7882), .D(n29818), 
         .Z(n13957)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22359_2_lut_4_lut.init = 16'h1000;
    LUT4 i5_2_lut_4_lut (.A(n31512), .B(clk_255kHz), .C(n7882), .D(n29530), 
         .Z(n14)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i5_2_lut_4_lut.init = 16'h0010;
    LUT4 i22485_2_lut_4_lut (.A(n31512), .B(clk_255kHz), .C(n7882), .D(n29944), 
         .Z(n14500)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22485_2_lut_4_lut.init = 16'h1000;
    CCU2D add_19627_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27125), .COUT(n27126));
    defparam add_19627_22.INIT0 = 16'h5555;
    defparam add_19627_22.INIT1 = 16'h5555;
    defparam add_19627_22.INJECT1_0 = "NO";
    defparam add_19627_22.INJECT1_1 = "NO";
    CCU2D add_19627_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27124), .COUT(n27125));
    defparam add_19627_20.INIT0 = 16'h5555;
    defparam add_19627_20.INIT1 = 16'h5555;
    defparam add_19627_20.INJECT1_0 = "NO";
    defparam add_19627_20.INJECT1_1 = "NO";
    CCU2D add_19627_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27123), .COUT(n27124));
    defparam add_19627_18.INIT0 = 16'h5555;
    defparam add_19627_18.INIT1 = 16'h5555;
    defparam add_19627_18.INJECT1_0 = "NO";
    defparam add_19627_18.INJECT1_1 = "NO";
    CCU2D add_19627_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27122), .COUT(n27123));
    defparam add_19627_16.INIT0 = 16'h5555;
    defparam add_19627_16.INIT1 = 16'h5555;
    defparam add_19627_16.INJECT1_0 = "NO";
    defparam add_19627_16.INJECT1_1 = "NO";
    CCU2D add_19627_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27121), .COUT(n27122));
    defparam add_19627_14.INIT0 = 16'h5555;
    defparam add_19627_14.INIT1 = 16'h5555;
    defparam add_19627_14.INJECT1_0 = "NO";
    defparam add_19627_14.INJECT1_1 = "NO";
    CCU2D add_19627_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27120), .COUT(n27121));
    defparam add_19627_12.INIT0 = 16'h5555;
    defparam add_19627_12.INIT1 = 16'h5555;
    defparam add_19627_12.INJECT1_0 = "NO";
    defparam add_19627_12.INJECT1_1 = "NO";
    CCU2D add_19627_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27119), .COUT(n27120));
    defparam add_19627_10.INIT0 = 16'h5555;
    defparam add_19627_10.INIT1 = 16'h5555;
    defparam add_19627_10.INJECT1_0 = "NO";
    defparam add_19627_10.INJECT1_1 = "NO";
    CCU2D add_19627_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27118), 
          .COUT(n27119));
    defparam add_19627_8.INIT0 = 16'h5555;
    defparam add_19627_8.INIT1 = 16'h5555;
    defparam add_19627_8.INJECT1_0 = "NO";
    defparam add_19627_8.INJECT1_1 = "NO";
    CCU2D add_19627_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27117), 
          .COUT(n27118));
    defparam add_19627_6.INIT0 = 16'h5555;
    defparam add_19627_6.INIT1 = 16'h5555;
    defparam add_19627_6.INJECT1_0 = "NO";
    defparam add_19627_6.INJECT1_1 = "NO";
    CCU2D add_19627_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27116), 
          .COUT(n27117));
    defparam add_19627_4.INIT0 = 16'h5555;
    defparam add_19627_4.INIT1 = 16'h5aaa;
    defparam add_19627_4.INJECT1_0 = "NO";
    defparam add_19627_4.INJECT1_1 = "NO";
    CCU2D add_19627_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27116));
    defparam add_19627_2.INIT0 = 16'h7000;
    defparam add_19627_2.INIT1 = 16'h5aaa;
    defparam add_19627_2.INJECT1_0 = "NO";
    defparam add_19627_2.INJECT1_1 = "NO";
    LUT4 i22325_2_lut_4_lut (.A(n31512), .B(clk_255kHz), .C(n7882), .D(n29784), 
         .Z(n27564)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22325_2_lut_4_lut.init = 16'h1000;
    LUT4 i22352_2_lut_4_lut (.A(n31512), .B(clk_255kHz), .C(n7882), .D(n29811), 
         .Z(n27547)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22352_2_lut_4_lut.init = 16'h1000;
    CCU2D count_2671_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26907), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_33.INIT1 = 16'h0000;
    defparam count_2671_add_4_33.INJECT1_0 = "NO";
    defparam count_2671_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26906), .COUT(n26907), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_31.INJECT1_0 = "NO";
    defparam count_2671_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26905), .COUT(n26906), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_29.INJECT1_0 = "NO";
    defparam count_2671_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26904), .COUT(n26905), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_27.INJECT1_0 = "NO";
    defparam count_2671_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26903), .COUT(n26904), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_25.INJECT1_0 = "NO";
    defparam count_2671_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26902), .COUT(n26903), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_23.INJECT1_0 = "NO";
    defparam count_2671_add_4_23.INJECT1_1 = "NO";
    FD1S3IX count_2671__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2824), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i1.GSR = "ENABLED";
    FD1S3IX count_2671__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2824), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i2.GSR = "ENABLED";
    FD1S3IX count_2671__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2824), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i3.GSR = "ENABLED";
    FD1S3IX count_2671__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2824), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i4.GSR = "ENABLED";
    FD1S3IX count_2671__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2824), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i5.GSR = "ENABLED";
    FD1S3IX count_2671__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2824), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i6.GSR = "ENABLED";
    FD1S3IX count_2671__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2824), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i7.GSR = "ENABLED";
    FD1S3IX count_2671__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2824), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i8.GSR = "ENABLED";
    FD1S3IX count_2671__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2824), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i9.GSR = "ENABLED";
    FD1S3IX count_2671__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i10.GSR = "ENABLED";
    FD1S3IX count_2671__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i11.GSR = "ENABLED";
    FD1S3IX count_2671__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i12.GSR = "ENABLED";
    FD1S3IX count_2671__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i13.GSR = "ENABLED";
    FD1S3IX count_2671__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i14.GSR = "ENABLED";
    FD1S3IX count_2671__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i15.GSR = "ENABLED";
    FD1S3IX count_2671__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i16.GSR = "ENABLED";
    FD1S3IX count_2671__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i17.GSR = "ENABLED";
    FD1S3IX count_2671__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i18.GSR = "ENABLED";
    FD1S3IX count_2671__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i19.GSR = "ENABLED";
    FD1S3IX count_2671__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i20.GSR = "ENABLED";
    FD1S3IX count_2671__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i21.GSR = "ENABLED";
    FD1S3IX count_2671__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i22.GSR = "ENABLED";
    FD1S3IX count_2671__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i23.GSR = "ENABLED";
    FD1S3IX count_2671__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i24.GSR = "ENABLED";
    FD1S3IX count_2671__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i25.GSR = "ENABLED";
    FD1S3IX count_2671__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i26.GSR = "ENABLED";
    FD1S3IX count_2671__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i27.GSR = "ENABLED";
    FD1S3IX count_2671__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i28.GSR = "ENABLED";
    FD1S3IX count_2671__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i29.GSR = "ENABLED";
    FD1S3IX count_2671__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i30.GSR = "ENABLED";
    FD1S3IX count_2671__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2824), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671__i31.GSR = "ENABLED";
    CCU2D count_2671_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26901), .COUT(n26902), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_21.INJECT1_0 = "NO";
    defparam count_2671_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26900), .COUT(n26901), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_19.INJECT1_0 = "NO";
    defparam count_2671_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26899), .COUT(n26900), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_17.INJECT1_0 = "NO";
    defparam count_2671_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26898), .COUT(n26899), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_15.INJECT1_0 = "NO";
    defparam count_2671_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26897), .COUT(n26898), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_13.INJECT1_0 = "NO";
    defparam count_2671_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26896), .COUT(n26897), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_11.INJECT1_0 = "NO";
    defparam count_2671_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26895), .COUT(n26896), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_9.INJECT1_0 = "NO";
    defparam count_2671_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26894), .COUT(n26895), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_7.INJECT1_0 = "NO";
    defparam count_2671_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26893), .COUT(n26894), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_5.INJECT1_0 = "NO";
    defparam count_2671_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26892), .COUT(n26893), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2671_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2671_add_4_3.INJECT1_0 = "NO";
    defparam count_2671_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2671_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26892), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2671_add_4_1.INIT0 = 16'hF000;
    defparam count_2671_add_4_1.INIT1 = 16'h0555;
    defparam count_2671_add_4_1.INJECT1_0 = "NO";
    defparam count_2671_add_4_1.INJECT1_1 = "NO";
    LUT4 i22368_2_lut_4_lut (.A(n31512), .B(clk_255kHz), .C(n7882), .D(n29827), 
         .Z(n27543)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22368_2_lut_4_lut.init = 16'h1000;
    LUT4 i22379_2_lut_4_lut (.A(n31512), .B(clk_255kHz), .C(n7882), .D(n29838), 
         .Z(n27550)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i22379_2_lut_4_lut.init = 16'h1000;
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0) 
//

module \ArmPeripheral(axis_haddr=8'b0)  (debug_c_c, n31512, databus, n4181, 
            \read_size[0] , n13941, n9379, Stepper_X_M0_c_0, n13917, 
            prev_step_clk, step_clk, limit_latched, prev_limit_latched, 
            n9297, prev_select, n31474, \register_addr[1] , Stepper_X_Dir_c, 
            \register_addr[0] , n1, Stepper_X_En_c, Stepper_X_M1_c_1, 
            \control_reg[7] , n12159, Stepper_X_M2_c_2, \read_size[2] , 
            n31435, n34, n27445, n29137, limit_c_0, read_value, 
            n31425, n24, n31421, VCC_net, GND_net, Stepper_X_nFault_c, 
            Stepper_X_Step_c, n31409, n8056, n8090, n17035) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n31512;
    input [31:0]databus;
    input n4181;
    output \read_size[0] ;
    input n13941;
    input n9379;
    output Stepper_X_M0_c_0;
    input n13917;
    output prev_step_clk;
    output step_clk;
    output limit_latched;
    output prev_limit_latched;
    input n9297;
    output prev_select;
    input n31474;
    input \register_addr[1] ;
    output Stepper_X_Dir_c;
    input \register_addr[0] ;
    input n1;
    output Stepper_X_En_c;
    output Stepper_X_M1_c_1;
    output \control_reg[7] ;
    input n12159;
    output Stepper_X_M2_c_2;
    output \read_size[2] ;
    input n31435;
    input n34;
    output n27445;
    input n29137;
    input limit_c_0;
    output [31:0]read_value;
    input n31425;
    input n24;
    input n31421;
    input VCC_net;
    input GND_net;
    input Stepper_X_nFault_c;
    output Stepper_X_Step_c;
    input n31409;
    output n8056;
    output n8090;
    input n17035;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n4182;
    wire [31:0]n224;
    
    wire n182;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n1_c, n2;
    wire [31:0]n6499;
    
    wire n29696, n29697, n1_adj_22, n2_adj_23, n2_adj_25;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n1_adj_26, n29684, n29685, n29686, n2_adj_27, fault_latched, 
        n29765, n29766, n49, n62, n58, n50, n41, n60, n54, 
        n42, n52, n38, n56, n46, n29698, n1_adj_28, n2_adj_29, 
        n29767, n29142, n29144, n29145, n29147, n29143, n29148, 
        n29149, n29151, n29146, n29152, n29150, n29153, n29154, 
        n29155, n29156, n29140, n29138, n29141, n29158, n29159, 
        n29160, n29161, n29139, n29157, int_step, n26883, n26882, 
        n26881, n26880, n26879, n26878, n26877, n26876, n26875, 
        n26874, n26873, n26872, n26871, n26870, n26869, n26868;
    
    FD1S3IX steps_reg__i26 (.D(n4182[26]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n4182[25]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n4182[24]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n4182[23]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n4182[22]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n4182[21]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n4182[20]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n4182[19]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n4182[18]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n4182[17]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n4182[16]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n4182[15]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n4182[14]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n4182[13]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n4182[12]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n4182[11]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n4182[10]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n4182[9]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n4182[8]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n4182[7]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n4182[6]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n4182[5]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n4182[4]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n4182[3]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n4182[2]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n4182[1]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 mux_1622_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n4181), .Z(n4182[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i10_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i0 (.D(n4182[0]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n9379), .SP(n13941), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3IX control_reg_i1 (.D(databus[0]), .SP(n13917), .CD(n31512), 
            .CK(debug_c_c), .Q(Stepper_X_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i0 (.D(databus[0]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n31474), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    LUT4 mux_1622_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n4181), .Z(n4182[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i9_3_lut.init = 16'hcaca;
    PFUMX mux_1930_Mux_5_i3 (.BLUT(n1_c), .ALUT(n2), .C0(\register_addr[1] ), 
          .Z(n6499[5]));
    LUT4 i22136_3_lut (.A(Stepper_X_M0_c_0), .B(div_factor_reg[0]), .C(\register_addr[1] ), 
         .Z(n29696)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22136_3_lut.init = 16'hcaca;
    LUT4 i22137_3_lut (.A(limit_latched), .B(steps_reg[0]), .C(\register_addr[1] ), 
         .Z(n29697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22137_3_lut.init = 16'hcaca;
    LUT4 i15139_2_lut (.A(Stepper_X_Dir_c), .B(\register_addr[0] ), .Z(n1_c)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15139_2_lut.init = 16'h2222;
    LUT4 mux_1930_Mux_5_i2_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), 
         .C(\register_addr[0] ), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1930_Mux_5_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n4181), .Z(n4182[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i8_3_lut.init = 16'hcaca;
    PFUMX mux_1930_Mux_6_i3 (.BLUT(n1_adj_22), .ALUT(n2_adj_23), .C0(\register_addr[1] ), 
          .Z(n6499[6]));
    LUT4 mux_1622_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n4181), .Z(n4182[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i7_3_lut.init = 16'hcaca;
    PFUMX mux_1930_Mux_7_i3 (.BLUT(n1), .ALUT(n2_adj_25), .C0(\register_addr[1] ), 
          .Z(n6499[7]));
    LUT4 mux_1622_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n4181), 
         .Z(n4182[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n4181), .Z(n4182[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n4181), .Z(n4182[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n4181), 
         .Z(n4182[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n4181), 
         .Z(n4182[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n4181), .Z(n4182[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n4181), 
         .Z(n4182[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n4181), .Z(n4182[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n4181), .Z(n4182[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n4181), 
         .Z(n4182[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n4181), 
         .Z(n4182[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n4181), 
         .Z(n4182[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n4181), 
         .Z(n4182[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i13_3_lut.init = 16'hcaca;
    LUT4 i15136_2_lut (.A(Stepper_X_En_c), .B(\register_addr[0] ), .Z(n1_adj_22)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15136_2_lut.init = 16'h2222;
    LUT4 mux_1930_Mux_6_i2_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), 
         .C(\register_addr[0] ), .Z(n2_adj_23)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1930_Mux_6_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1930_Mux_7_i2_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), 
         .C(\register_addr[0] ), .Z(n2_adj_25)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1930_Mux_7_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n4181), 
         .Z(n4182[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n4181), 
         .Z(n4182[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i11_3_lut.init = 16'hcaca;
    LUT4 i15141_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n1_adj_26)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15141_2_lut.init = 16'h2222;
    PFUMX i22126 (.BLUT(n29684), .ALUT(n29685), .C0(\register_addr[1] ), 
          .Z(n29686));
    LUT4 mux_1930_Mux_3_i2_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), 
         .C(\register_addr[0] ), .Z(n2_adj_27)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1930_Mux_3_i2_3_lut.init = 16'hcaca;
    LUT4 i22205_3_lut (.A(Stepper_X_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n29765)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22205_3_lut.init = 16'hcaca;
    LUT4 i22206_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n29766)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22206_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n4181), 
         .Z(n4182[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n4181), 
         .Z(n4182[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i17_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n9297), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n9297), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n9297), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n9297), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n9297), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n9297), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n9297), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n9297), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n13917), .CD(n12159), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n13917), .PD(n31512), 
            .CK(debug_c_c), .Q(Stepper_X_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n13917), .PD(n31512), 
            .CK(debug_c_c), .Q(Stepper_X_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n13917), .CD(n31512), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n13917), .PD(n31512), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n13917), .CD(n31512), 
            .CK(debug_c_c), .Q(Stepper_X_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n13917), .PD(n31512), 
            .CK(debug_c_c), .Q(Stepper_X_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n31435), .SP(n13941), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    LUT4 mux_1622_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n4181), 
         .Z(n4182[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i21_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i31 (.D(n4182[31]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n4182[30]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n4182[29]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n4182[28]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    LUT4 i22124_3_lut (.A(Stepper_X_M2_c_2), .B(n34), .C(\register_addr[0] ), 
         .Z(n29684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22124_3_lut.init = 16'hcaca;
    LUT4 i22125_3_lut (.A(div_factor_reg[2]), .B(steps_reg[2]), .C(\register_addr[0] ), 
         .Z(n29685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22125_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n27445)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 mux_1622_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n4181), 
         .Z(n4182[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n4181), 
         .Z(n4182[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n4181), 
         .Z(n4182[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i29_3_lut.init = 16'hcaca;
    LUT4 i17_4_lut (.A(steps_reg[8]), .B(steps_reg[27]), .C(steps_reg[31]), 
         .D(steps_reg[30]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[15]), .B(n52), .C(n38), .D(steps_reg[11]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[20]), .B(steps_reg[18]), .C(steps_reg[24]), 
         .D(steps_reg[4]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[9]), .B(steps_reg[12]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[5]), .B(n56), .C(n46), .D(steps_reg[6]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[7]), .B(steps_reg[26]), .C(steps_reg[25]), 
         .D(steps_reg[16]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[17]), .B(steps_reg[21]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    PFUMX i22138 (.BLUT(n29696), .ALUT(n29697), .C0(\register_addr[0] ), 
          .Z(n29698));
    LUT4 mux_1622_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n4181), 
         .Z(n4182[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i15_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i27 (.D(n4182[27]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    LUT4 i24_4_lut (.A(steps_reg[19]), .B(steps_reg[3]), .C(steps_reg[22]), 
         .D(steps_reg[13]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[10]), .B(steps_reg[14]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[29]), .B(steps_reg[0]), .C(steps_reg[2]), 
         .D(steps_reg[1]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[28]), .B(steps_reg[23]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 mux_1622_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n4181), .Z(n4182[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i1_3_lut.init = 16'hcaca;
    LUT4 i15140_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n1_adj_28)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15140_2_lut.init = 16'h2222;
    LUT4 mux_1930_Mux_4_i2_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), 
         .C(\register_addr[0] ), .Z(n2_adj_29)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1930_Mux_4_i2_3_lut.init = 16'hcaca;
    PFUMX mux_1930_Mux_3_i3 (.BLUT(n1_adj_26), .ALUT(n2_adj_27), .C0(\register_addr[1] ), 
          .Z(n6499[3]));
    PFUMX i22207 (.BLUT(n29765), .ALUT(n29766), .C0(\register_addr[1] ), 
          .Z(n29767));
    LUT4 i1_4_lut (.A(div_factor_reg[31]), .B(n29137), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n29142)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'hc088;
    LUT4 mux_1622_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n4181), 
         .Z(n4182[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i20_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_32 (.A(div_factor_reg[30]), .B(n29137), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n29144)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_32.init = 16'hc088;
    LUT4 i1_4_lut_adj_33 (.A(div_factor_reg[29]), .B(n29137), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n29145)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_33.init = 16'hc088;
    LUT4 i1_4_lut_adj_34 (.A(div_factor_reg[28]), .B(n29137), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n29147)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_34.init = 16'hc088;
    LUT4 i118_1_lut (.A(limit_c_0), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_35 (.A(div_factor_reg[27]), .B(n29137), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n29143)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_35.init = 16'hc088;
    FD1P3AX read_value__i31 (.D(n29142), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n29144), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n29145), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n29147), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n29143), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n29148), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n29149), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29151), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29146), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29152), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29150), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29153), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    LUT4 mux_1622_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n4181), 
         .Z(n4182[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i16_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i19 (.D(n29154), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29155), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29156), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29140), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29138), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29141), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29158), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29159), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29160), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29161), .SP(n13941), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29139), .SP(n13941), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29157), .SP(n13941), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6499[7]), .SP(n13941), .CD(n31425), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6499[6]), .SP(n13941), .CD(n31425), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n6499[5]), .SP(n13941), .CD(n31425), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6499[4]), .SP(n13941), .CD(n31425), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6499[3]), .SP(n13941), .CD(n31425), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n29686), .SP(n13941), .CD(n31425), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n29767), .SP(n13941), .CD(n31425), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_36 (.A(div_factor_reg[26]), .B(n29137), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n29148)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_36.init = 16'hc088;
    FD1P3AX int_step_182 (.D(n31421), .SP(n24), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_X_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_37 (.A(div_factor_reg[25]), .B(n29137), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n29149)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_37.init = 16'hc088;
    LUT4 i1_4_lut_adj_38 (.A(div_factor_reg[24]), .B(n29137), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n29151)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_38.init = 16'hc088;
    LUT4 i1_4_lut_adj_39 (.A(div_factor_reg[23]), .B(n29137), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n29146)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_39.init = 16'hc088;
    LUT4 i1_4_lut_adj_40 (.A(div_factor_reg[22]), .B(n29137), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n29152)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_40.init = 16'hc088;
    LUT4 i1_4_lut_adj_41 (.A(div_factor_reg[21]), .B(n29137), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n29150)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_41.init = 16'hc088;
    LUT4 i1_4_lut_adj_42 (.A(div_factor_reg[20]), .B(n29137), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n29153)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_42.init = 16'hc088;
    LUT4 i1_4_lut_adj_43 (.A(div_factor_reg[19]), .B(n29137), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n29154)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_43.init = 16'hc088;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26883), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_44 (.A(div_factor_reg[18]), .B(n29137), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n29155)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_44.init = 16'hc088;
    LUT4 i1_4_lut_adj_45 (.A(div_factor_reg[17]), .B(n29137), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n29156)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_45.init = 16'hc088;
    LUT4 i1_4_lut_adj_46 (.A(div_factor_reg[16]), .B(n29137), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n29140)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_4_lut_adj_46.init = 16'hc088;
    LUT4 i1_4_lut_adj_47 (.A(div_factor_reg[15]), .B(n29137), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n29138)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_47.init = 16'hc088;
    LUT4 i1_4_lut_adj_48 (.A(div_factor_reg[14]), .B(n29137), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n29141)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_48.init = 16'hc088;
    LUT4 i1_4_lut_adj_49 (.A(div_factor_reg[13]), .B(n29137), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n29158)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_49.init = 16'hc088;
    LUT4 i1_4_lut_adj_50 (.A(div_factor_reg[12]), .B(n29137), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n29159)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_50.init = 16'hc088;
    LUT4 i1_4_lut_adj_51 (.A(div_factor_reg[11]), .B(n29137), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n29160)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_51.init = 16'hc088;
    LUT4 i1_4_lut_adj_52 (.A(div_factor_reg[10]), .B(n29137), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n29161)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_52.init = 16'hc088;
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26882), .COUT(n26883), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_53 (.A(div_factor_reg[9]), .B(n29137), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n29139)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_53.init = 16'hc088;
    LUT4 i1_4_lut_adj_54 (.A(div_factor_reg[8]), .B(n29137), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n29157)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_54.init = 16'hc088;
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26881), .COUT(n26882), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26880), .COUT(n26881), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26879), .COUT(n26880), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26878), .COUT(n26879), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    FD1P3IX read_value__i0 (.D(n29698), .SP(n13941), .CD(n31425), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26877), .COUT(n26878), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26876), .COUT(n26877), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26875), .COUT(n26876), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26874), .COUT(n26875), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26873), .COUT(n26874), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26872), .COUT(n26873), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26871), .COUT(n26872), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26870), .COUT(n26871), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26869), .COUT(n26870), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    LUT4 mux_1622_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n4181), 
         .Z(n4182[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i19_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26868), .COUT(n26869), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(step_clk), .C1(n34), .D1(prev_step_clk), 
          .COUT(n26868), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    PFUMX mux_1930_Mux_4_i3 (.BLUT(n1_adj_28), .ALUT(n2_adj_29), .C0(\register_addr[1] ), 
          .Z(n6499[4]));
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_X_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 mux_1622_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n4181), 
         .Z(n4182[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1622_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n4181), 
         .Z(n4182[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1622_i25_3_lut.init = 16'hcaca;
    ClockDivider_U8 step_clk_gen (.GND_net(GND_net), .step_clk(step_clk), 
            .debug_c_c(debug_c_c), .n31512(n31512), .n31409(n31409), .n8056(n8056), 
            .div_factor_reg({div_factor_reg}), .n8090(n8090), .n17035(n17035)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U8
//

module ClockDivider_U8 (GND_net, step_clk, debug_c_c, n31512, n31409, 
            n8056, div_factor_reg, n8090, n17035) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output step_clk;
    input debug_c_c;
    input n31512;
    input n31409;
    output n8056;
    input [31:0]div_factor_reg;
    output n8090;
    input n17035;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26996;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n26997, n26995, n26994, n26993, n26992, n26991, n26990, 
        n26989, n26988, n8021, n26819;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    wire [31:0]n40;
    
    wire n26818, n26699, n26817, n26698, n26697, n26696, n26816, 
        n26815, n26814, n26813, n26812, n26811, n26695, n26694, 
        n26810, n26809, n26693, n26808, n26807, n26806, n26692, 
        n26805, n26691, n26804, n26690, n26689, n26688, n26687, 
        n26686, n26685, n26684, n26683, n26682, n26681, n26680, 
        n26679, n26678, n26677, n26676, n26675, n26674, n26673, 
        n26672, n26671, n26670, n26669, n26668, n26667, n26666, 
        n26665, n26664, n26663, n26662, n26661, n26660, n26659, 
        n26658, n26657, n26656, n26655, n26654, n26653, n26652, 
        n27003, n27002, n27001, n27000, n26999, n26998;
    
    CCU2D count_2674_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26996), .COUT(n26997), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_19.INJECT1_0 = "NO";
    defparam count_2674_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26995), .COUT(n26996), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_17.INJECT1_0 = "NO";
    defparam count_2674_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26994), .COUT(n26995), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_15.INJECT1_0 = "NO";
    defparam count_2674_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26993), .COUT(n26994), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_13.INJECT1_0 = "NO";
    defparam count_2674_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26992), .COUT(n26993), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_11.INJECT1_0 = "NO";
    defparam count_2674_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26991), .COUT(n26992), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_9.INJECT1_0 = "NO";
    defparam count_2674_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26990), .COUT(n26991), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_7.INJECT1_0 = "NO";
    defparam count_2674_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26989), .COUT(n26990), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_5.INJECT1_0 = "NO";
    defparam count_2674_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26988), .COUT(n26989), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_3.INJECT1_0 = "NO";
    defparam count_2674_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26988), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_1.INIT0 = 16'hF000;
    defparam count_2674_add_4_1.INIT1 = 16'h0555;
    defparam count_2674_add_4_1.INJECT1_0 = "NO";
    defparam count_2674_add_4_1.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n8021), .CK(debug_c_c), .CD(n31512), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26819), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26818), .COUT(n26819), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26699), .S1(n8021));
    defparam sub_2064_add_2_33.INIT0 = 16'h5555;
    defparam sub_2064_add_2_33.INIT1 = 16'h0000;
    defparam sub_2064_add_2_33.INJECT1_0 = "NO";
    defparam sub_2064_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26817), .COUT(n26818), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26698), .COUT(n26699));
    defparam sub_2064_add_2_31.INIT0 = 16'h5999;
    defparam sub_2064_add_2_31.INIT1 = 16'h5999;
    defparam sub_2064_add_2_31.INJECT1_0 = "NO";
    defparam sub_2064_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26697), .COUT(n26698));
    defparam sub_2064_add_2_29.INIT0 = 16'h5999;
    defparam sub_2064_add_2_29.INIT1 = 16'h5999;
    defparam sub_2064_add_2_29.INJECT1_0 = "NO";
    defparam sub_2064_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26696), .COUT(n26697));
    defparam sub_2064_add_2_27.INIT0 = 16'h5999;
    defparam sub_2064_add_2_27.INIT1 = 16'h5999;
    defparam sub_2064_add_2_27.INJECT1_0 = "NO";
    defparam sub_2064_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26816), .COUT(n26817), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26815), .COUT(n26816), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26814), .COUT(n26815), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26813), .COUT(n26814), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26812), .COUT(n26813), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26811), .COUT(n26812), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26695), .COUT(n26696));
    defparam sub_2064_add_2_25.INIT0 = 16'h5999;
    defparam sub_2064_add_2_25.INIT1 = 16'h5999;
    defparam sub_2064_add_2_25.INJECT1_0 = "NO";
    defparam sub_2064_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26694), .COUT(n26695));
    defparam sub_2064_add_2_23.INIT0 = 16'h5999;
    defparam sub_2064_add_2_23.INIT1 = 16'h5999;
    defparam sub_2064_add_2_23.INJECT1_0 = "NO";
    defparam sub_2064_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26810), .COUT(n26811), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26809), .COUT(n26810), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26693), .COUT(n26694));
    defparam sub_2064_add_2_21.INIT0 = 16'h5999;
    defparam sub_2064_add_2_21.INIT1 = 16'h5999;
    defparam sub_2064_add_2_21.INJECT1_0 = "NO";
    defparam sub_2064_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26808), .COUT(n26809), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26807), .COUT(n26808), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26806), .COUT(n26807), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26692), .COUT(n26693));
    defparam sub_2064_add_2_19.INIT0 = 16'h5999;
    defparam sub_2064_add_2_19.INIT1 = 16'h5999;
    defparam sub_2064_add_2_19.INJECT1_0 = "NO";
    defparam sub_2064_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26805), .COUT(n26806), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26691), .COUT(n26692));
    defparam sub_2064_add_2_17.INIT0 = 16'h5999;
    defparam sub_2064_add_2_17.INIT1 = 16'h5999;
    defparam sub_2064_add_2_17.INJECT1_0 = "NO";
    defparam sub_2064_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26804), .COUT(n26805), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26804), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26690), .COUT(n26691));
    defparam sub_2064_add_2_15.INIT0 = 16'h5999;
    defparam sub_2064_add_2_15.INIT1 = 16'h5999;
    defparam sub_2064_add_2_15.INJECT1_0 = "NO";
    defparam sub_2064_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26689), .COUT(n26690));
    defparam sub_2064_add_2_13.INIT0 = 16'h5999;
    defparam sub_2064_add_2_13.INIT1 = 16'h5999;
    defparam sub_2064_add_2_13.INJECT1_0 = "NO";
    defparam sub_2064_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26688), .COUT(n26689));
    defparam sub_2064_add_2_11.INIT0 = 16'h5999;
    defparam sub_2064_add_2_11.INIT1 = 16'h5999;
    defparam sub_2064_add_2_11.INJECT1_0 = "NO";
    defparam sub_2064_add_2_11.INJECT1_1 = "NO";
    FD1S3IX count_2674__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i0.GSR = "ENABLED";
    CCU2D sub_2064_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26687), .COUT(n26688));
    defparam sub_2064_add_2_9.INIT0 = 16'h5999;
    defparam sub_2064_add_2_9.INIT1 = 16'h5999;
    defparam sub_2064_add_2_9.INJECT1_0 = "NO";
    defparam sub_2064_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26686), .COUT(n26687));
    defparam sub_2064_add_2_7.INIT0 = 16'h5999;
    defparam sub_2064_add_2_7.INIT1 = 16'h5999;
    defparam sub_2064_add_2_7.INJECT1_0 = "NO";
    defparam sub_2064_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26685), .COUT(n26686));
    defparam sub_2064_add_2_5.INIT0 = 16'h5999;
    defparam sub_2064_add_2_5.INIT1 = 16'h5999;
    defparam sub_2064_add_2_5.INJECT1_0 = "NO";
    defparam sub_2064_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26684), .COUT(n26685));
    defparam sub_2064_add_2_3.INIT0 = 16'h5999;
    defparam sub_2064_add_2_3.INIT1 = 16'h5999;
    defparam sub_2064_add_2_3.INJECT1_0 = "NO";
    defparam sub_2064_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26684));
    defparam sub_2064_add_2_1.INIT0 = 16'h0000;
    defparam sub_2064_add_2_1.INIT1 = 16'h5999;
    defparam sub_2064_add_2_1.INJECT1_0 = "NO";
    defparam sub_2064_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26683), .S1(n8056));
    defparam sub_2066_add_2_33.INIT0 = 16'h5999;
    defparam sub_2066_add_2_33.INIT1 = 16'h0000;
    defparam sub_2066_add_2_33.INJECT1_0 = "NO";
    defparam sub_2066_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26682), .COUT(n26683));
    defparam sub_2066_add_2_31.INIT0 = 16'h5999;
    defparam sub_2066_add_2_31.INIT1 = 16'h5999;
    defparam sub_2066_add_2_31.INJECT1_0 = "NO";
    defparam sub_2066_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26681), .COUT(n26682));
    defparam sub_2066_add_2_29.INIT0 = 16'h5999;
    defparam sub_2066_add_2_29.INIT1 = 16'h5999;
    defparam sub_2066_add_2_29.INJECT1_0 = "NO";
    defparam sub_2066_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26680), .COUT(n26681));
    defparam sub_2066_add_2_27.INIT0 = 16'h5999;
    defparam sub_2066_add_2_27.INIT1 = 16'h5999;
    defparam sub_2066_add_2_27.INJECT1_0 = "NO";
    defparam sub_2066_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26679), .COUT(n26680));
    defparam sub_2066_add_2_25.INIT0 = 16'h5999;
    defparam sub_2066_add_2_25.INIT1 = 16'h5999;
    defparam sub_2066_add_2_25.INJECT1_0 = "NO";
    defparam sub_2066_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26678), .COUT(n26679));
    defparam sub_2066_add_2_23.INIT0 = 16'h5999;
    defparam sub_2066_add_2_23.INIT1 = 16'h5999;
    defparam sub_2066_add_2_23.INJECT1_0 = "NO";
    defparam sub_2066_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26677), .COUT(n26678));
    defparam sub_2066_add_2_21.INIT0 = 16'h5999;
    defparam sub_2066_add_2_21.INIT1 = 16'h5999;
    defparam sub_2066_add_2_21.INJECT1_0 = "NO";
    defparam sub_2066_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26676), .COUT(n26677));
    defparam sub_2066_add_2_19.INIT0 = 16'h5999;
    defparam sub_2066_add_2_19.INIT1 = 16'h5999;
    defparam sub_2066_add_2_19.INJECT1_0 = "NO";
    defparam sub_2066_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26675), .COUT(n26676));
    defparam sub_2066_add_2_17.INIT0 = 16'h5999;
    defparam sub_2066_add_2_17.INIT1 = 16'h5999;
    defparam sub_2066_add_2_17.INJECT1_0 = "NO";
    defparam sub_2066_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26674), .COUT(n26675));
    defparam sub_2066_add_2_15.INIT0 = 16'h5999;
    defparam sub_2066_add_2_15.INIT1 = 16'h5999;
    defparam sub_2066_add_2_15.INJECT1_0 = "NO";
    defparam sub_2066_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26673), .COUT(n26674));
    defparam sub_2066_add_2_13.INIT0 = 16'h5999;
    defparam sub_2066_add_2_13.INIT1 = 16'h5999;
    defparam sub_2066_add_2_13.INJECT1_0 = "NO";
    defparam sub_2066_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26672), .COUT(n26673));
    defparam sub_2066_add_2_11.INIT0 = 16'h5999;
    defparam sub_2066_add_2_11.INIT1 = 16'h5999;
    defparam sub_2066_add_2_11.INJECT1_0 = "NO";
    defparam sub_2066_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26671), .COUT(n26672));
    defparam sub_2066_add_2_9.INIT0 = 16'h5999;
    defparam sub_2066_add_2_9.INIT1 = 16'h5999;
    defparam sub_2066_add_2_9.INJECT1_0 = "NO";
    defparam sub_2066_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26670), .COUT(n26671));
    defparam sub_2066_add_2_7.INIT0 = 16'h5999;
    defparam sub_2066_add_2_7.INIT1 = 16'h5999;
    defparam sub_2066_add_2_7.INJECT1_0 = "NO";
    defparam sub_2066_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26669), .COUT(n26670));
    defparam sub_2066_add_2_5.INIT0 = 16'h5999;
    defparam sub_2066_add_2_5.INIT1 = 16'h5999;
    defparam sub_2066_add_2_5.INJECT1_0 = "NO";
    defparam sub_2066_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26668), .COUT(n26669));
    defparam sub_2066_add_2_3.INIT0 = 16'h5999;
    defparam sub_2066_add_2_3.INIT1 = 16'h5999;
    defparam sub_2066_add_2_3.INJECT1_0 = "NO";
    defparam sub_2066_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2066_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n26668));
    defparam sub_2066_add_2_1.INIT0 = 16'h0000;
    defparam sub_2066_add_2_1.INIT1 = 16'h5999;
    defparam sub_2066_add_2_1.INJECT1_0 = "NO";
    defparam sub_2066_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26667), .S1(n8090));
    defparam sub_2067_add_2_33.INIT0 = 16'hf555;
    defparam sub_2067_add_2_33.INIT1 = 16'h0000;
    defparam sub_2067_add_2_33.INJECT1_0 = "NO";
    defparam sub_2067_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26666), .COUT(n26667));
    defparam sub_2067_add_2_31.INIT0 = 16'hf555;
    defparam sub_2067_add_2_31.INIT1 = 16'hf555;
    defparam sub_2067_add_2_31.INJECT1_0 = "NO";
    defparam sub_2067_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26665), .COUT(n26666));
    defparam sub_2067_add_2_29.INIT0 = 16'hf555;
    defparam sub_2067_add_2_29.INIT1 = 16'hf555;
    defparam sub_2067_add_2_29.INJECT1_0 = "NO";
    defparam sub_2067_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26664), .COUT(n26665));
    defparam sub_2067_add_2_27.INIT0 = 16'hf555;
    defparam sub_2067_add_2_27.INIT1 = 16'hf555;
    defparam sub_2067_add_2_27.INJECT1_0 = "NO";
    defparam sub_2067_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26663), .COUT(n26664));
    defparam sub_2067_add_2_25.INIT0 = 16'hf555;
    defparam sub_2067_add_2_25.INIT1 = 16'hf555;
    defparam sub_2067_add_2_25.INJECT1_0 = "NO";
    defparam sub_2067_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26662), .COUT(n26663));
    defparam sub_2067_add_2_23.INIT0 = 16'hf555;
    defparam sub_2067_add_2_23.INIT1 = 16'hf555;
    defparam sub_2067_add_2_23.INJECT1_0 = "NO";
    defparam sub_2067_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26661), .COUT(n26662));
    defparam sub_2067_add_2_21.INIT0 = 16'hf555;
    defparam sub_2067_add_2_21.INIT1 = 16'hf555;
    defparam sub_2067_add_2_21.INJECT1_0 = "NO";
    defparam sub_2067_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26660), .COUT(n26661));
    defparam sub_2067_add_2_19.INIT0 = 16'hf555;
    defparam sub_2067_add_2_19.INIT1 = 16'hf555;
    defparam sub_2067_add_2_19.INJECT1_0 = "NO";
    defparam sub_2067_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26659), .COUT(n26660));
    defparam sub_2067_add_2_17.INIT0 = 16'hf555;
    defparam sub_2067_add_2_17.INIT1 = 16'hf555;
    defparam sub_2067_add_2_17.INJECT1_0 = "NO";
    defparam sub_2067_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26658), .COUT(n26659));
    defparam sub_2067_add_2_15.INIT0 = 16'hf555;
    defparam sub_2067_add_2_15.INIT1 = 16'hf555;
    defparam sub_2067_add_2_15.INJECT1_0 = "NO";
    defparam sub_2067_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26657), .COUT(n26658));
    defparam sub_2067_add_2_13.INIT0 = 16'hf555;
    defparam sub_2067_add_2_13.INIT1 = 16'hf555;
    defparam sub_2067_add_2_13.INJECT1_0 = "NO";
    defparam sub_2067_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26656), .COUT(n26657));
    defparam sub_2067_add_2_11.INIT0 = 16'hf555;
    defparam sub_2067_add_2_11.INIT1 = 16'hf555;
    defparam sub_2067_add_2_11.INJECT1_0 = "NO";
    defparam sub_2067_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26655), .COUT(n26656));
    defparam sub_2067_add_2_9.INIT0 = 16'hf555;
    defparam sub_2067_add_2_9.INIT1 = 16'hf555;
    defparam sub_2067_add_2_9.INJECT1_0 = "NO";
    defparam sub_2067_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26654), .COUT(n26655));
    defparam sub_2067_add_2_7.INIT0 = 16'hf555;
    defparam sub_2067_add_2_7.INIT1 = 16'hf555;
    defparam sub_2067_add_2_7.INJECT1_0 = "NO";
    defparam sub_2067_add_2_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    CCU2D sub_2067_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26653), .COUT(n26654));
    defparam sub_2067_add_2_5.INIT0 = 16'hf555;
    defparam sub_2067_add_2_5.INIT1 = 16'hf555;
    defparam sub_2067_add_2_5.INJECT1_0 = "NO";
    defparam sub_2067_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26652), .COUT(n26653));
    defparam sub_2067_add_2_3.INIT0 = 16'hf555;
    defparam sub_2067_add_2_3.INIT1 = 16'hf555;
    defparam sub_2067_add_2_3.INJECT1_0 = "NO";
    defparam sub_2067_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n26652));
    defparam sub_2067_add_2_1.INIT0 = 16'h0000;
    defparam sub_2067_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2067_add_2_1.INJECT1_0 = "NO";
    defparam sub_2067_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31409), .PD(n17035), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    FD1S3IX count_2674__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i1.GSR = "ENABLED";
    FD1S3IX count_2674__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i2.GSR = "ENABLED";
    FD1S3IX count_2674__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i3.GSR = "ENABLED";
    FD1S3IX count_2674__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i4.GSR = "ENABLED";
    FD1S3IX count_2674__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i5.GSR = "ENABLED";
    FD1S3IX count_2674__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i6.GSR = "ENABLED";
    FD1S3IX count_2674__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i7.GSR = "ENABLED";
    FD1S3IX count_2674__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i8.GSR = "ENABLED";
    FD1S3IX count_2674__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i9.GSR = "ENABLED";
    FD1S3IX count_2674__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i10.GSR = "ENABLED";
    FD1S3IX count_2674__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i11.GSR = "ENABLED";
    FD1S3IX count_2674__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i12.GSR = "ENABLED";
    FD1S3IX count_2674__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i13.GSR = "ENABLED";
    FD1S3IX count_2674__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i14.GSR = "ENABLED";
    FD1S3IX count_2674__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i15.GSR = "ENABLED";
    FD1S3IX count_2674__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i16.GSR = "ENABLED";
    FD1S3IX count_2674__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i17.GSR = "ENABLED";
    FD1S3IX count_2674__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i18.GSR = "ENABLED";
    FD1S3IX count_2674__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i19.GSR = "ENABLED";
    FD1S3IX count_2674__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i20.GSR = "ENABLED";
    FD1S3IX count_2674__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i21.GSR = "ENABLED";
    FD1S3IX count_2674__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i22.GSR = "ENABLED";
    FD1S3IX count_2674__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i23.GSR = "ENABLED";
    FD1S3IX count_2674__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i24.GSR = "ENABLED";
    FD1S3IX count_2674__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i25.GSR = "ENABLED";
    FD1S3IX count_2674__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i26.GSR = "ENABLED";
    FD1S3IX count_2674__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i27.GSR = "ENABLED";
    FD1S3IX count_2674__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i28.GSR = "ENABLED";
    FD1S3IX count_2674__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i29.GSR = "ENABLED";
    FD1S3IX count_2674__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i30.GSR = "ENABLED";
    FD1S3IX count_2674__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31409), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674__i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31409), .CD(n17035), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D count_2674_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27003), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_33.INIT1 = 16'h0000;
    defparam count_2674_add_4_33.INJECT1_0 = "NO";
    defparam count_2674_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27002), .COUT(n27003), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_31.INJECT1_0 = "NO";
    defparam count_2674_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27001), .COUT(n27002), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_29.INJECT1_0 = "NO";
    defparam count_2674_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27000), .COUT(n27001), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_27.INJECT1_0 = "NO";
    defparam count_2674_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26999), .COUT(n27000), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_25.INJECT1_0 = "NO";
    defparam count_2674_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26998), .COUT(n26999), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_23.INJECT1_0 = "NO";
    defparam count_2674_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2674_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26997), .COUT(n26998), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2674_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2674_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2674_add_4_21.INJECT1_0 = "NO";
    defparam count_2674_add_4_21.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module EncoderPeripheral
//

module EncoderPeripheral (\register_addr[0] , n31432, prev_select, debug_c_c, 
            n31471, \read_size[0] , n15087, n6, encoder_rb_c, encoder_ra_c, 
            read_value, \read_size[2] , n31541, encoder_ri_c, qreset, 
            VCC_net, GND_net, \quadA_delayed[1] , n13939, n6_adj_4, 
            \quadB_delayed[1] ) /* synthesis syn_module_defined=1 */ ;
    input \register_addr[0] ;
    input n31432;
    output prev_select;
    input debug_c_c;
    input n31471;
    output \read_size[0] ;
    input n15087;
    input n6;
    input encoder_rb_c;
    input encoder_ra_c;
    output [31:0]read_value;
    output \read_size[2] ;
    input n31541;
    input encoder_ri_c;
    input qreset;
    input VCC_net;
    input GND_net;
    output \quadA_delayed[1] ;
    input n13939;
    output n6_adj_4;
    output \quadB_delayed[1] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(58[14:22])
    
    wire n29086, n29081, n29106, n29103, n29092, n29085, n29089, 
        n29095, n29105, n29082, n29093, n29094, n29096, n29097, 
        n29083, n29084, n29091, n29099, n29107, n29100, n29087, 
        n29108, n29090, n29109, n29101, n29098, n29088, n29102, 
        n29104;
    wire [31:0]n180;
    
    LUT4 i1_2_lut_3_lut (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [4]), 
         .Z(n29086)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_4 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [5]), 
         .Z(n29081)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_4.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_5 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [6]), 
         .Z(n29106)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_5.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_6 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [7]), 
         .Z(n29103)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_6.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_7 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [8]), 
         .Z(n29092)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_7.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_8 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [9]), 
         .Z(n29085)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_8.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_9 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [10]), 
         .Z(n29089)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_9.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_10 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [11]), 
         .Z(n29095)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_10.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_11 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [12]), 
         .Z(n29105)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_11.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_12 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [13]), 
         .Z(n29082)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_12.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_13 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [14]), 
         .Z(n29093)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_13.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_14 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [15]), 
         .Z(n29094)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_14.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_15 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [16]), 
         .Z(n29096)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_15.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_16 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [17]), 
         .Z(n29097)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_16.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_17 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [18]), 
         .Z(n29083)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_17.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_18 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [19]), 
         .Z(n29084)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_18.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_19 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [20]), 
         .Z(n29091)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_19.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_20 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [21]), 
         .Z(n29099)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_20.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_21 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [22]), 
         .Z(n29107)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_21.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_22 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [23]), 
         .Z(n29100)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_22.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_23 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [24]), 
         .Z(n29087)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_23.init = 16'h2020;
    FD1S3AX prev_select_126 (.D(n31471), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam prev_select_126.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_24 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [25]), 
         .Z(n29108)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_24.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_25 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [26]), 
         .Z(n29090)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_25.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_26 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [27]), 
         .Z(n29109)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_26.init = 16'h2020;
    FD1P3IX read_size__i1 (.D(n6), .SP(n15087), .CD(n31432), .CK(debug_c_c), 
            .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_size__i1.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_27 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [28]), 
         .Z(n29101)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_27.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_28 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [29]), 
         .Z(n29098)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_28.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_29 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [30]), 
         .Z(n29088)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_29.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_30 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [31]), 
         .Z(n29102)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_30.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_31 (.A(\register_addr[0] ), .B(n31432), .C(\register[1] [0]), 
         .Z(n29104)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_31.init = 16'h2020;
    LUT4 mux_115_Mux_2_i1_3_lut (.A(encoder_rb_c), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n180[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_3_i1_3_lut (.A(encoder_ra_c), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n180[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_3_i1_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i1 (.D(n180[1]), .SP(n15087), .CD(n31432), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_size__i2 (.D(n31541), .SP(n15087), .CD(n31432), .CK(debug_c_c), 
            .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n180[2]), .SP(n15087), .CD(n31432), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n180[3]), .SP(n15087), .CD(n31432), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3AX read_value__i4 (.D(n29086), .SP(n15087), .CK(debug_c_c), .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3AX read_value__i5 (.D(n29081), .SP(n15087), .CK(debug_c_c), .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3AX read_value__i6 (.D(n29106), .SP(n15087), .CK(debug_c_c), .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3AX read_value__i7 (.D(n29103), .SP(n15087), .CK(debug_c_c), .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29092), .SP(n15087), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29085), .SP(n15087), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29089), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29095), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29105), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29082), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29093), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29094), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29096), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29097), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29083), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n29084), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29091), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29099), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29107), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29100), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29087), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n29108), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n29090), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n29109), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n29101), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n29098), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n29088), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n29102), .SP(n15087), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX read_value__i0 (.D(n29104), .SP(n15087), .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 mux_115_Mux_1_i1_3_lut (.A(encoder_ri_c), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n180[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_1_i1_3_lut.init = 16'hcaca;
    QuadratureDecoder q (.\register[1] ({\register[1] }), .debug_c_c(debug_c_c), 
            .qreset(qreset), .VCC_net(VCC_net), .GND_net(GND_net), .encoder_rb_c(encoder_rb_c), 
            .encoder_ra_c(encoder_ra_c), .\quadA_delayed[1] (\quadA_delayed[1] ), 
            .n13939(n13939), .n6(n6_adj_4), .\quadB_delayed[1] (\quadB_delayed[1] )) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(92[20] 96[37])
    
endmodule
//
// Verilog Description of module QuadratureDecoder
//

module QuadratureDecoder (\register[1] , debug_c_c, qreset, VCC_net, 
            GND_net, encoder_rb_c, encoder_ra_c, \quadA_delayed[1] , 
            n13939, n6, \quadB_delayed[1] ) /* synthesis syn_module_defined=1 */ ;
    output [31:0]\register[1] ;
    input debug_c_c;
    input qreset;
    input VCC_net;
    input GND_net;
    input encoder_rb_c;
    input encoder_ra_c;
    output \quadA_delayed[1] ;
    input n13939;
    output n6;
    output \quadB_delayed[1] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(15[13:18])
    wire [2:0]quadB_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    wire [2:0]quadA_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    
    wire n26522;
    wire [31:0]n4424;
    
    wire n26521, n26520, n26519, n26518, n26517, n26516, n26515, 
        n26514, n26513, n26512, n26511, n26510, n26509, n26508, 
        n26507;
    
    FD1P3AX count_at_reset_i0_i0 (.D(count[0]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i0.GSR = "ENABLED";
    IFS1P3DX quadB_delayed_i0 (.D(encoder_rb_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadB_delayed[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i0.GSR = "ENABLED";
    IFS1P3DX quadA_delayed_i0 (.D(encoder_ra_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadA_delayed[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i0.GSR = "ENABLED";
    CCU2D add_1718_33 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[30]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[31]), .D1(GND_net), .CIN(n26522), .S0(n4424[30]), 
          .S1(n4424[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_33.INIT0 = 16'h6969;
    defparam add_1718_33.INIT1 = 16'h6969;
    defparam add_1718_33.INJECT1_0 = "NO";
    defparam add_1718_33.INJECT1_1 = "NO";
    CCU2D add_1718_31 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[28]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[29]), .D1(GND_net), .CIN(n26521), .COUT(n26522), 
          .S0(n4424[28]), .S1(n4424[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_31.INIT0 = 16'h6969;
    defparam add_1718_31.INIT1 = 16'h6969;
    defparam add_1718_31.INJECT1_0 = "NO";
    defparam add_1718_31.INJECT1_1 = "NO";
    CCU2D add_1718_29 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[26]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[27]), .D1(GND_net), .CIN(n26520), .COUT(n26521), 
          .S0(n4424[26]), .S1(n4424[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_29.INIT0 = 16'h6969;
    defparam add_1718_29.INIT1 = 16'h6969;
    defparam add_1718_29.INJECT1_0 = "NO";
    defparam add_1718_29.INJECT1_1 = "NO";
    CCU2D add_1718_27 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[24]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[25]), .D1(GND_net), .CIN(n26519), .COUT(n26520), 
          .S0(n4424[24]), .S1(n4424[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_27.INIT0 = 16'h6969;
    defparam add_1718_27.INIT1 = 16'h6969;
    defparam add_1718_27.INJECT1_0 = "NO";
    defparam add_1718_27.INJECT1_1 = "NO";
    CCU2D add_1718_25 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[22]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[23]), .D1(GND_net), .CIN(n26518), .COUT(n26519), 
          .S0(n4424[22]), .S1(n4424[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_25.INIT0 = 16'h6969;
    defparam add_1718_25.INIT1 = 16'h6969;
    defparam add_1718_25.INJECT1_0 = "NO";
    defparam add_1718_25.INJECT1_1 = "NO";
    CCU2D add_1718_23 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[20]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[21]), .D1(GND_net), .CIN(n26517), .COUT(n26518), 
          .S0(n4424[20]), .S1(n4424[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_23.INIT0 = 16'h6969;
    defparam add_1718_23.INIT1 = 16'h6969;
    defparam add_1718_23.INJECT1_0 = "NO";
    defparam add_1718_23.INJECT1_1 = "NO";
    CCU2D add_1718_21 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[18]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[19]), .D1(GND_net), .CIN(n26516), .COUT(n26517), 
          .S0(n4424[18]), .S1(n4424[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_21.INIT0 = 16'h6969;
    defparam add_1718_21.INIT1 = 16'h6969;
    defparam add_1718_21.INJECT1_0 = "NO";
    defparam add_1718_21.INJECT1_1 = "NO";
    CCU2D add_1718_19 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[16]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[17]), .D1(GND_net), .CIN(n26515), .COUT(n26516), 
          .S0(n4424[16]), .S1(n4424[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_19.INIT0 = 16'h6969;
    defparam add_1718_19.INIT1 = 16'h6969;
    defparam add_1718_19.INJECT1_0 = "NO";
    defparam add_1718_19.INJECT1_1 = "NO";
    CCU2D add_1718_17 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[14]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[15]), .D1(GND_net), .CIN(n26514), .COUT(n26515), 
          .S0(n4424[14]), .S1(n4424[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_17.INIT0 = 16'h6969;
    defparam add_1718_17.INIT1 = 16'h6969;
    defparam add_1718_17.INJECT1_0 = "NO";
    defparam add_1718_17.INJECT1_1 = "NO";
    CCU2D add_1718_15 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[12]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[13]), .D1(GND_net), .CIN(n26513), .COUT(n26514), 
          .S0(n4424[12]), .S1(n4424[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_15.INIT0 = 16'h6969;
    defparam add_1718_15.INIT1 = 16'h6969;
    defparam add_1718_15.INJECT1_0 = "NO";
    defparam add_1718_15.INJECT1_1 = "NO";
    CCU2D add_1718_13 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[10]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[11]), .D1(GND_net), .CIN(n26512), .COUT(n26513), 
          .S0(n4424[10]), .S1(n4424[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_13.INIT0 = 16'h6969;
    defparam add_1718_13.INIT1 = 16'h6969;
    defparam add_1718_13.INJECT1_0 = "NO";
    defparam add_1718_13.INJECT1_1 = "NO";
    CCU2D add_1718_11 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[8]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[9]), .D1(GND_net), .CIN(n26511), .COUT(n26512), 
          .S0(n4424[8]), .S1(n4424[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_11.INIT0 = 16'h6969;
    defparam add_1718_11.INIT1 = 16'h6969;
    defparam add_1718_11.INJECT1_0 = "NO";
    defparam add_1718_11.INJECT1_1 = "NO";
    CCU2D add_1718_9 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[6]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[7]), .D1(GND_net), .CIN(n26510), .COUT(n26511), 
          .S0(n4424[6]), .S1(n4424[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_9.INIT0 = 16'h6969;
    defparam add_1718_9.INIT1 = 16'h6969;
    defparam add_1718_9.INJECT1_0 = "NO";
    defparam add_1718_9.INJECT1_1 = "NO";
    CCU2D add_1718_7 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[4]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[5]), .D1(GND_net), .CIN(n26509), .COUT(n26510), 
          .S0(n4424[4]), .S1(n4424[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_7.INIT0 = 16'h6969;
    defparam add_1718_7.INIT1 = 16'h6969;
    defparam add_1718_7.INJECT1_0 = "NO";
    defparam add_1718_7.INJECT1_1 = "NO";
    CCU2D add_1718_5 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[2]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[3]), .D1(GND_net), .CIN(n26508), .COUT(n26509), 
          .S0(n4424[2]), .S1(n4424[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_5.INIT0 = 16'h6969;
    defparam add_1718_5.INIT1 = 16'h6969;
    defparam add_1718_5.INJECT1_0 = "NO";
    defparam add_1718_5.INJECT1_1 = "NO";
    CCU2D add_1718_3 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[0]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[1]), .D1(GND_net), .CIN(n26507), .COUT(n26508), 
          .S0(n4424[0]), .S1(n4424[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_3.INIT0 = 16'h9696;
    defparam add_1718_3.INIT1 = 16'h6969;
    defparam add_1718_3.INJECT1_0 = "NO";
    defparam add_1718_3.INJECT1_1 = "NO";
    CCU2D add_1718_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26507));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1718_1.INIT0 = 16'hF000;
    defparam add_1718_1.INIT1 = 16'h6666;
    defparam add_1718_1.INJECT1_0 = "NO";
    defparam add_1718_1.INJECT1_1 = "NO";
    FD1P3IX count__i31 (.D(n4424[31]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i31.GSR = "ENABLED";
    FD1P3IX count__i30 (.D(n4424[30]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i30.GSR = "ENABLED";
    FD1P3IX count__i29 (.D(n4424[29]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i29.GSR = "ENABLED";
    FD1P3IX count__i28 (.D(n4424[28]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i28.GSR = "ENABLED";
    FD1P3IX count__i27 (.D(n4424[27]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i27.GSR = "ENABLED";
    FD1P3IX count__i26 (.D(n4424[26]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i26.GSR = "ENABLED";
    FD1P3IX count__i25 (.D(n4424[25]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i25.GSR = "ENABLED";
    FD1P3IX count__i24 (.D(n4424[24]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i24.GSR = "ENABLED";
    FD1P3IX count__i23 (.D(n4424[23]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i23.GSR = "ENABLED";
    FD1P3IX count__i22 (.D(n4424[22]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i22.GSR = "ENABLED";
    FD1P3IX count__i21 (.D(n4424[21]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i21.GSR = "ENABLED";
    FD1P3IX count__i20 (.D(n4424[20]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i20.GSR = "ENABLED";
    FD1P3IX count__i19 (.D(n4424[19]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i19.GSR = "ENABLED";
    FD1P3IX count__i18 (.D(n4424[18]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i18.GSR = "ENABLED";
    FD1P3IX count__i17 (.D(n4424[17]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i17.GSR = "ENABLED";
    FD1P3IX count__i16 (.D(n4424[16]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i16.GSR = "ENABLED";
    FD1P3IX count__i15 (.D(n4424[15]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i15.GSR = "ENABLED";
    FD1P3IX count__i14 (.D(n4424[14]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i14.GSR = "ENABLED";
    FD1P3IX count__i13 (.D(n4424[13]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i13.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n4424[12]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i12.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n4424[11]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n4424[10]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n4424[9]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n4424[8]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n4424[7]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n4424[6]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n4424[5]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n4424[4]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n4424[3]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n4424[2]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n4424[1]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i1.GSR = "ENABLED";
    LUT4 i2_2_lut (.A(quadB_delayed[2]), .B(quadA_delayed[2]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(18[22:95])
    defparam i2_2_lut.init = 16'h6666;
    FD1P3IX count__i0 (.D(n4424[0]), .SP(n13939), .CD(qreset), .CK(debug_c_c), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i0.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i1 (.D(count[1]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i1.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i2 (.D(count[2]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i2.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i3 (.D(count[3]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i3.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i4 (.D(count[4]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i4.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i5 (.D(count[5]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i5.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i6 (.D(count[6]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i6.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i7 (.D(count[7]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i7.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i8 (.D(count[8]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i8.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i9 (.D(count[9]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i9.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i10 (.D(count[10]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i10.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i11 (.D(count[11]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i11.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i12 (.D(count[12]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i12.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i13 (.D(count[13]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i13.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i14 (.D(count[14]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i14.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i15 (.D(count[15]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i15.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i16 (.D(count[16]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i16.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i17 (.D(count[17]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i17.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i18 (.D(count[18]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i18.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i19 (.D(count[19]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i19.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i20 (.D(count[20]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i20.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i21 (.D(count[21]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i21.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i22 (.D(count[22]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i22.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i23 (.D(count[23]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i23.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i24 (.D(count[24]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i24.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i25 (.D(count[25]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i25.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i26 (.D(count[26]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i26.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i27 (.D(count[27]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i27.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i28 (.D(count[28]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i28.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i29 (.D(count[29]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i29.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i30 (.D(count[30]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i30.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i31 (.D(count[31]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i31.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i1 (.D(quadB_delayed[0]), .CK(debug_c_c), .Q(\quadB_delayed[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i2 (.D(\quadB_delayed[1] ), .CK(debug_c_c), .Q(quadB_delayed[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i2.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i1 (.D(quadA_delayed[0]), .CK(debug_c_c), .Q(\quadA_delayed[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i2 (.D(\quadA_delayed[1] ), .CK(debug_c_c), .Q(quadA_delayed[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i2.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ClockDividerP_SP(factor=120000) 
//

module \ClockDividerP_SP(factor=120000)  (n29792, debug_c_0, debug_c_c, 
            n31512, n2861, GND_net) /* synthesis syn_module_defined=1 */ ;
    output n29792;
    output debug_c_0;
    input debug_c_c;
    input n31512;
    input n2861;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(86[13:18])
    
    wire n21, n19, n25, n38, n34, n26, n31481, n20, n36, n30, 
        n32, n22, n29536, n29680, n29534, n29662, n29542, n27789;
    wire [31:0]n134;
    
    wire n26939, n26938, n26937, n26936, n26935, n26934, n26933, 
        n26932, n26931, n26930, n26929, n26928, n26927, n26926, 
        n26925, n26924;
    
    LUT4 i9_4_lut (.A(count[5]), .B(count[16]), .C(count[12]), .D(count[14]), 
         .Z(n21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i7_4_lut (.A(count[7]), .B(count[15]), .C(count[4]), .D(count[10]), 
         .Z(n19)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut_rep_337 (.A(n25), .B(n38), .C(n34), .D(n26), .Z(n31481)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i19_4_lut_rep_337.init = 16'hfffe;
    LUT4 i8_4_lut (.A(count[1]), .B(count[0]), .C(count[2]), .D(count[3]), 
         .Z(n20)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(count[11]), .B(count[13]), .Z(n25)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i18_4_lut (.A(count[6]), .B(n36), .C(n30), .D(count[9]), .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(count[20]), .B(count[31]), .C(count[24]), .D(count[30]), 
         .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(count[21]), .B(count[17]), .Z(n26)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i16_4_lut (.A(count[26]), .B(n32), .C(n22), .D(count[29]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(count[18]), .B(count[28]), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i12_4_lut (.A(count[25]), .B(count[23]), .C(count[8]), .D(count[27]), 
         .Z(n32)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[19]), .B(count[22]), .Z(n22)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(102[9:26])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i22332_4_lut (.A(n31481), .B(n29536), .C(n29680), .D(n29534), 
         .Z(n29792)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i22332_4_lut.init = 16'h4000;
    LUT4 i21982_2_lut (.A(count[10]), .B(count[12]), .Z(n29536)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21982_2_lut.init = 16'h8888;
    LUT4 i22120_4_lut (.A(count[3]), .B(n29662), .C(n29542), .D(count[0]), 
         .Z(n29680)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22120_4_lut.init = 16'h8000;
    LUT4 i21980_2_lut (.A(count[2]), .B(count[5]), .Z(n29534)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21980_2_lut.init = 16'h8888;
    LUT4 i22102_4_lut (.A(count[1]), .B(count[16]), .C(count[4]), .D(count[15]), 
         .Z(n29662)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22102_4_lut.init = 16'h8000;
    LUT4 i21988_2_lut (.A(count[7]), .B(count[14]), .Z(n29542)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21988_2_lut.init = 16'h8888;
    FD1S3IX clk_o_13 (.D(n27789), .CK(debug_c_c), .CD(n31512), .Q(debug_c_0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(88[9] 107[6])
    defparam clk_o_13.GSR = "ENABLED";
    FD1S3IX count_2672__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2861), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i0.GSR = "ENABLED";
    CCU2D count_2672_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26939), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_33.INIT1 = 16'h0000;
    defparam count_2672_add_4_33.INJECT1_0 = "NO";
    defparam count_2672_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26938), .COUT(n26939), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_31.INJECT1_0 = "NO";
    defparam count_2672_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26937), .COUT(n26938), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_29.INJECT1_0 = "NO";
    defparam count_2672_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26936), .COUT(n26937), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_27.INJECT1_0 = "NO";
    defparam count_2672_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26935), .COUT(n26936), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_25.INJECT1_0 = "NO";
    defparam count_2672_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26934), .COUT(n26935), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_23.INJECT1_0 = "NO";
    defparam count_2672_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26933), .COUT(n26934), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_21.INJECT1_0 = "NO";
    defparam count_2672_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26932), .COUT(n26933), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_19.INJECT1_0 = "NO";
    defparam count_2672_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26931), .COUT(n26932), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_17.INJECT1_0 = "NO";
    defparam count_2672_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26930), .COUT(n26931), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_15.INJECT1_0 = "NO";
    defparam count_2672_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26929), .COUT(n26930), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_13.INJECT1_0 = "NO";
    defparam count_2672_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26928), .COUT(n26929), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_11.INJECT1_0 = "NO";
    defparam count_2672_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26927), .COUT(n26928), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_9.INJECT1_0 = "NO";
    defparam count_2672_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26926), .COUT(n26927), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_7.INJECT1_0 = "NO";
    defparam count_2672_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26925), .COUT(n26926), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_5.INJECT1_0 = "NO";
    defparam count_2672_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26924), .COUT(n26925), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2672_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2672_add_4_3.INJECT1_0 = "NO";
    defparam count_2672_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2672_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26924), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672_add_4_1.INIT0 = 16'hF000;
    defparam count_2672_add_4_1.INIT1 = 16'h0555;
    defparam count_2672_add_4_1.INJECT1_0 = "NO";
    defparam count_2672_add_4_1.INJECT1_1 = "NO";
    LUT4 i22376_4_lut_4_lut (.A(n31481), .B(n20), .C(n19), .D(n21), 
         .Z(n27789)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i22376_4_lut_4_lut.init = 16'h0001;
    FD1S3IX count_2672__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2861), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i1.GSR = "ENABLED";
    FD1S3IX count_2672__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2861), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i2.GSR = "ENABLED";
    FD1S3IX count_2672__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2861), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i3.GSR = "ENABLED";
    FD1S3IX count_2672__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2861), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i4.GSR = "ENABLED";
    FD1S3IX count_2672__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2861), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i5.GSR = "ENABLED";
    FD1S3IX count_2672__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2861), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i6.GSR = "ENABLED";
    FD1S3IX count_2672__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2861), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i7.GSR = "ENABLED";
    FD1S3IX count_2672__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2861), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i8.GSR = "ENABLED";
    FD1S3IX count_2672__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2861), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i9.GSR = "ENABLED";
    FD1S3IX count_2672__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i10.GSR = "ENABLED";
    FD1S3IX count_2672__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i11.GSR = "ENABLED";
    FD1S3IX count_2672__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i12.GSR = "ENABLED";
    FD1S3IX count_2672__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i13.GSR = "ENABLED";
    FD1S3IX count_2672__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i14.GSR = "ENABLED";
    FD1S3IX count_2672__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i15.GSR = "ENABLED";
    FD1S3IX count_2672__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i16.GSR = "ENABLED";
    FD1S3IX count_2672__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i17.GSR = "ENABLED";
    FD1S3IX count_2672__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i18.GSR = "ENABLED";
    FD1S3IX count_2672__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i19.GSR = "ENABLED";
    FD1S3IX count_2672__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i20.GSR = "ENABLED";
    FD1S3IX count_2672__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i21.GSR = "ENABLED";
    FD1S3IX count_2672__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i22.GSR = "ENABLED";
    FD1S3IX count_2672__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i23.GSR = "ENABLED";
    FD1S3IX count_2672__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i24.GSR = "ENABLED";
    FD1S3IX count_2672__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i25.GSR = "ENABLED";
    FD1S3IX count_2672__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i26.GSR = "ENABLED";
    FD1S3IX count_2672__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i27.GSR = "ENABLED";
    FD1S3IX count_2672__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i28.GSR = "ENABLED";
    FD1S3IX count_2672__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i29.GSR = "ENABLED";
    FD1S3IX count_2672__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i30.GSR = "ENABLED";
    FD1S3IX count_2672__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2861), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2672__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module EncoderPeripheral_U11
//

module EncoderPeripheral_U11 (\read_size[0] , debug_c_c, n14146, n31427, 
            n31450, prev_select, n31465, \read_size[2] , n31478, read_value, 
            \register_addr[0] , encoder_la_c, encoder_lb_c, n59, n57, 
            n45, \quadA_delayed[1] , qreset, n6, \quadB_delayed[1] , 
            n13939, n97, encoder_li_c, GND_net, \register[1][0] , 
            VCC_net, \register[1][19] , \register[1][20] , \register[1][26] ) /* synthesis syn_module_defined=1 */ ;
    output \read_size[0] ;
    input debug_c_c;
    input n14146;
    input n31427;
    input n31450;
    output prev_select;
    input n31465;
    output \read_size[2] ;
    input n31478;
    output [31:0]read_value;
    input \register_addr[0] ;
    input encoder_la_c;
    input encoder_lb_c;
    input n59;
    input n57;
    input n45;
    input \quadA_delayed[1] ;
    input qreset;
    input n6;
    input \quadB_delayed[1] ;
    output n13939;
    input n97;
    input encoder_li_c;
    input GND_net;
    output \register[1][0] ;
    input VCC_net;
    output \register[1][19] ;
    output \register[1][20] ;
    output \register[1][26] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]n100;
    wire [31:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(58[14:22])
    wire [2:0]quadA_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    
    wire n6_adj_19;
    wire [2:0]quadB_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    
    wire n15145;
    
    FD1P3IX read_size__i1 (.D(n31450), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1S3AX prev_select_126 (.D(n31465), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam prev_select_126.GSR = "ENABLED";
    FD1P3IX read_size__i2 (.D(n31478), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i28.GSR = "ENABLED";
    LUT4 i15002_2_lut (.A(\register[1] [31]), .B(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15002_2_lut.init = 16'h8888;
    LUT4 i15003_2_lut (.A(\register[1] [30]), .B(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15003_2_lut.init = 16'h8888;
    LUT4 i15004_2_lut (.A(\register[1] [29]), .B(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15004_2_lut.init = 16'h8888;
    LUT4 i15007_2_lut (.A(\register[1] [28]), .B(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15007_2_lut.init = 16'h8888;
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n100[23]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n100[7]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n100[2]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n100[1]), .SP(n14146), .CD(n31427), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i15008_2_lut (.A(\register[1] [27]), .B(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15008_2_lut.init = 16'h8888;
    LUT4 i15009_2_lut (.A(\register[1] [25]), .B(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15009_2_lut.init = 16'h8888;
    LUT4 i15010_2_lut (.A(\register[1] [24]), .B(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15010_2_lut.init = 16'h8888;
    LUT4 i15011_2_lut (.A(\register[1] [23]), .B(\register_addr[0] ), .Z(n100[23])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15011_2_lut.init = 16'h8888;
    LUT4 i15012_2_lut (.A(\register[1] [22]), .B(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15012_2_lut.init = 16'h8888;
    LUT4 i15013_2_lut (.A(\register[1] [21]), .B(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15013_2_lut.init = 16'h8888;
    LUT4 i15014_2_lut (.A(\register[1] [18]), .B(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15014_2_lut.init = 16'h8888;
    LUT4 i15015_2_lut (.A(\register[1] [17]), .B(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15015_2_lut.init = 16'h8888;
    LUT4 i15016_2_lut (.A(\register[1] [16]), .B(\register_addr[0] ), .Z(n100[16])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15016_2_lut.init = 16'h8888;
    LUT4 i15017_2_lut (.A(\register[1] [15]), .B(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15017_2_lut.init = 16'h8888;
    LUT4 i15018_2_lut (.A(\register[1] [14]), .B(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15018_2_lut.init = 16'h8888;
    LUT4 i15019_2_lut (.A(\register[1] [13]), .B(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15019_2_lut.init = 16'h8888;
    LUT4 i15020_2_lut (.A(\register[1] [12]), .B(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15020_2_lut.init = 16'h8888;
    LUT4 i15021_2_lut (.A(\register[1] [11]), .B(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15021_2_lut.init = 16'h8888;
    LUT4 i15022_2_lut (.A(\register[1] [10]), .B(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15022_2_lut.init = 16'h8888;
    LUT4 i15023_2_lut (.A(\register[1] [9]), .B(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15023_2_lut.init = 16'h8888;
    LUT4 i15024_2_lut (.A(\register[1] [8]), .B(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15024_2_lut.init = 16'h8888;
    LUT4 i15025_2_lut (.A(\register[1] [7]), .B(\register_addr[0] ), .Z(n100[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15025_2_lut.init = 16'h8888;
    LUT4 i15026_2_lut (.A(\register[1] [6]), .B(\register_addr[0] ), .Z(n100[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15026_2_lut.init = 16'h8888;
    LUT4 i15027_2_lut (.A(\register[1] [5]), .B(\register_addr[0] ), .Z(n100[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15027_2_lut.init = 16'h8888;
    LUT4 i15028_2_lut (.A(\register[1] [4]), .B(\register_addr[0] ), .Z(n100[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15028_2_lut.init = 16'h8888;
    LUT4 mux_115_Mux_3_i1_3_lut (.A(encoder_la_c), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n100[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_2_i1_3_lut (.A(encoder_lb_c), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n100[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_2_i1_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i19 (.D(n59), .SP(n14146), .CK(debug_c_c), .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n57), .SP(n14146), .CK(debug_c_c), .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n45), .SP(n14146), .CK(debug_c_c), .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i26.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(\quadA_delayed[1] ), .B(qreset), .C(n6), .D(\quadB_delayed[1] ), 
         .Z(n13939)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(62[18:35])
    defparam i1_4_lut.init = 16'hedde;
    FD1P3AX read_value__i0 (.D(n97), .SP(n14146), .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 mux_115_Mux_1_i1_3_lut (.A(encoder_li_c), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n100[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_3 (.A(quadA_delayed[1]), .B(qreset), .C(n6_adj_19), 
         .D(quadB_delayed[1]), .Z(n15145)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(62[18:35])
    defparam i1_4_lut_adj_3.init = 16'hedde;
    QuadratureDecoder_U6 q (.GND_net(GND_net), .quadA_delayed({Open_2, quadA_delayed[1], 
            Open_3}), .\register[1] ({\register[1] [31:27], \register[1][26] , 
            \register[1] [25:21], \register[1][20] , \register[1][19] , 
            \register[1] [18:1], \register[1][0] }), .debug_c_c(debug_c_c), 
            .qreset(qreset), .VCC_net(VCC_net), .encoder_lb_c(encoder_lb_c), 
            .n15145(n15145), .encoder_la_c(encoder_la_c), .\quadB_delayed[1] (quadB_delayed[1]), 
            .n6(n6_adj_19)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(92[20] 96[37])
    
endmodule
//
// Verilog Description of module QuadratureDecoder_U6
//

module QuadratureDecoder_U6 (GND_net, quadA_delayed, \register[1] , debug_c_c, 
            qreset, VCC_net, encoder_lb_c, n15145, encoder_la_c, \quadB_delayed[1] , 
            n6) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output [2:0]quadA_delayed;
    output [31:0]\register[1] ;
    input debug_c_c;
    input qreset;
    input VCC_net;
    input encoder_lb_c;
    input n15145;
    input encoder_la_c;
    output \quadB_delayed[1] ;
    output n6;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [2:0]quadB_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    
    wire n26439;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(15[13:18])
    wire [31:0]n4358;
    wire [2:0]quadA_delayed_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    
    wire n26454, n26453;
    wire [31:0]n100;
    
    wire n26452, n26451, n26450, n26449, n26448, n26447, n26446, 
        n26445, n26444, n26443, n26442, n26441, n26440;
    
    CCU2D add_1684_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26439));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_1.INIT0 = 16'hF000;
    defparam add_1684_1.INIT1 = 16'h6666;
    defparam add_1684_1.INJECT1_0 = "NO";
    defparam add_1684_1.INJECT1_1 = "NO";
    FD1P3AX count_at_reset_i0_i0 (.D(count[0]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i0.GSR = "ENABLED";
    IFS1P3DX quadB_delayed_i0 (.D(encoder_lb_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadB_delayed[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i0.GSR = "ENABLED";
    FD1P3IX count__i0 (.D(n4358[0]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i0.GSR = "ENABLED";
    IFS1P3DX quadA_delayed_i0 (.D(encoder_la_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadA_delayed_c[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i0.GSR = "ENABLED";
    CCU2D add_1684_33 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[30]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[31]), .D1(GND_net), .CIN(n26454), .S0(n4358[30]), 
          .S1(n4358[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_33.INIT0 = 16'h6969;
    defparam add_1684_33.INIT1 = 16'h6969;
    defparam add_1684_33.INJECT1_0 = "NO";
    defparam add_1684_33.INJECT1_1 = "NO";
    CCU2D add_1684_31 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[28]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[29]), .D1(GND_net), .CIN(n26453), .COUT(n26454), 
          .S0(n100[28]), .S1(n100[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_31.INIT0 = 16'h6969;
    defparam add_1684_31.INIT1 = 16'h6969;
    defparam add_1684_31.INJECT1_0 = "NO";
    defparam add_1684_31.INJECT1_1 = "NO";
    CCU2D add_1684_29 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[26]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[27]), .D1(GND_net), .CIN(n26452), .COUT(n26453), 
          .S0(n100[26]), .S1(n100[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_29.INIT0 = 16'h6969;
    defparam add_1684_29.INIT1 = 16'h6969;
    defparam add_1684_29.INJECT1_0 = "NO";
    defparam add_1684_29.INJECT1_1 = "NO";
    CCU2D add_1684_27 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[24]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[25]), .D1(GND_net), .CIN(n26451), .COUT(n26452), 
          .S0(n100[24]), .S1(n100[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_27.INIT0 = 16'h6969;
    defparam add_1684_27.INIT1 = 16'h6969;
    defparam add_1684_27.INJECT1_0 = "NO";
    defparam add_1684_27.INJECT1_1 = "NO";
    CCU2D add_1684_25 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[22]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[23]), .D1(GND_net), .CIN(n26450), .COUT(n26451), 
          .S0(n100[22]), .S1(n100[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_25.INIT0 = 16'h6969;
    defparam add_1684_25.INIT1 = 16'h6969;
    defparam add_1684_25.INJECT1_0 = "NO";
    defparam add_1684_25.INJECT1_1 = "NO";
    FD1P3IX count__i31 (.D(n4358[31]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i31.GSR = "ENABLED";
    FD1P3IX count__i30 (.D(n4358[30]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i30.GSR = "ENABLED";
    CCU2D add_1684_23 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[20]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[21]), .D1(GND_net), .CIN(n26449), .COUT(n26450), 
          .S0(n100[20]), .S1(n100[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_23.INIT0 = 16'h6969;
    defparam add_1684_23.INIT1 = 16'h6969;
    defparam add_1684_23.INJECT1_0 = "NO";
    defparam add_1684_23.INJECT1_1 = "NO";
    CCU2D add_1684_21 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[18]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[19]), .D1(GND_net), .CIN(n26448), .COUT(n26449), 
          .S0(n100[18]), .S1(n100[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_21.INIT0 = 16'h6969;
    defparam add_1684_21.INIT1 = 16'h6969;
    defparam add_1684_21.INJECT1_0 = "NO";
    defparam add_1684_21.INJECT1_1 = "NO";
    CCU2D add_1684_19 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[16]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[17]), .D1(GND_net), .CIN(n26447), .COUT(n26448), 
          .S0(n100[16]), .S1(n100[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_19.INIT0 = 16'h6969;
    defparam add_1684_19.INIT1 = 16'h6969;
    defparam add_1684_19.INJECT1_0 = "NO";
    defparam add_1684_19.INJECT1_1 = "NO";
    CCU2D add_1684_17 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[14]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[15]), .D1(GND_net), .CIN(n26446), .COUT(n26447), 
          .S0(n100[14]), .S1(n100[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_17.INIT0 = 16'h6969;
    defparam add_1684_17.INIT1 = 16'h6969;
    defparam add_1684_17.INJECT1_0 = "NO";
    defparam add_1684_17.INJECT1_1 = "NO";
    CCU2D add_1684_15 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[12]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[13]), .D1(GND_net), .CIN(n26445), .COUT(n26446), 
          .S0(n100[12]), .S1(n100[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_15.INIT0 = 16'h6969;
    defparam add_1684_15.INIT1 = 16'h6969;
    defparam add_1684_15.INJECT1_0 = "NO";
    defparam add_1684_15.INJECT1_1 = "NO";
    CCU2D add_1684_13 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[10]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[11]), .D1(GND_net), .CIN(n26444), .COUT(n26445), 
          .S0(n100[10]), .S1(n100[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_13.INIT0 = 16'h6969;
    defparam add_1684_13.INIT1 = 16'h6969;
    defparam add_1684_13.INJECT1_0 = "NO";
    defparam add_1684_13.INJECT1_1 = "NO";
    CCU2D add_1684_11 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[8]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[9]), .D1(GND_net), .CIN(n26443), .COUT(n26444), 
          .S0(n100[8]), .S1(n100[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_11.INIT0 = 16'h6969;
    defparam add_1684_11.INIT1 = 16'h6969;
    defparam add_1684_11.INJECT1_0 = "NO";
    defparam add_1684_11.INJECT1_1 = "NO";
    CCU2D add_1684_9 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[6]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[7]), .D1(GND_net), .CIN(n26442), .COUT(n26443), 
          .S0(n100[6]), .S1(n100[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_9.INIT0 = 16'h6969;
    defparam add_1684_9.INIT1 = 16'h6969;
    defparam add_1684_9.INJECT1_0 = "NO";
    defparam add_1684_9.INJECT1_1 = "NO";
    CCU2D add_1684_7 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[4]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[5]), .D1(GND_net), .CIN(n26441), .COUT(n26442), 
          .S0(n100[4]), .S1(n100[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_7.INIT0 = 16'h6969;
    defparam add_1684_7.INIT1 = 16'h6969;
    defparam add_1684_7.INJECT1_0 = "NO";
    defparam add_1684_7.INJECT1_1 = "NO";
    FD1P3AX count_at_reset_i0_i1 (.D(count[1]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i1.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i2 (.D(count[2]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i2.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i3 (.D(count[3]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i3.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i4 (.D(count[4]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i4.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i5 (.D(count[5]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i5.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i6 (.D(count[6]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i6.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i7 (.D(count[7]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i7.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i8 (.D(count[8]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i8.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i9 (.D(count[9]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i9.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i10 (.D(count[10]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i10.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i11 (.D(count[11]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i11.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i12 (.D(count[12]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i12.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i13 (.D(count[13]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i13.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i14 (.D(count[14]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i14.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i15 (.D(count[15]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i15.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i16 (.D(count[16]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i16.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i17 (.D(count[17]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i17.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i18 (.D(count[18]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i18.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i19 (.D(count[19]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i19.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i20 (.D(count[20]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i20.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i21 (.D(count[21]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i21.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i22 (.D(count[22]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i22.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i23 (.D(count[23]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i23.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i24 (.D(count[24]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i24.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i25 (.D(count[25]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i25.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i26 (.D(count[26]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i26.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i27 (.D(count[27]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i27.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i28 (.D(count[28]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i28.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i29 (.D(count[29]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i29.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i30 (.D(count[30]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i30.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i31 (.D(count[31]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i31.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i1 (.D(quadB_delayed[0]), .CK(debug_c_c), .Q(\quadB_delayed[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i2 (.D(\quadB_delayed[1] ), .CK(debug_c_c), .Q(quadB_delayed[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i2.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n100[1]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i1.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n100[2]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n100[3]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n100[4]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n100[5]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n100[6]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n100[7]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n100[8]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n100[9]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n100[10]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n100[11]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n100[12]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i12.GSR = "ENABLED";
    FD1P3IX count__i13 (.D(n100[13]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i13.GSR = "ENABLED";
    FD1P3IX count__i14 (.D(n100[14]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i14.GSR = "ENABLED";
    FD1P3IX count__i15 (.D(n100[15]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i15.GSR = "ENABLED";
    FD1P3IX count__i16 (.D(n100[16]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i16.GSR = "ENABLED";
    FD1P3IX count__i17 (.D(n100[17]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i17.GSR = "ENABLED";
    FD1P3IX count__i18 (.D(n100[18]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i18.GSR = "ENABLED";
    FD1P3IX count__i19 (.D(n100[19]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i19.GSR = "ENABLED";
    FD1P3IX count__i20 (.D(n100[20]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i20.GSR = "ENABLED";
    FD1P3IX count__i21 (.D(n100[21]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i21.GSR = "ENABLED";
    FD1P3IX count__i22 (.D(n100[22]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i22.GSR = "ENABLED";
    FD1P3IX count__i23 (.D(n100[23]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i23.GSR = "ENABLED";
    FD1P3IX count__i24 (.D(n100[24]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i24.GSR = "ENABLED";
    FD1P3IX count__i25 (.D(n100[25]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i25.GSR = "ENABLED";
    FD1P3IX count__i26 (.D(n100[26]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i26.GSR = "ENABLED";
    FD1P3IX count__i27 (.D(n100[27]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i27.GSR = "ENABLED";
    FD1P3IX count__i28 (.D(n100[28]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i28.GSR = "ENABLED";
    FD1P3IX count__i29 (.D(n100[29]), .SP(n15145), .CD(qreset), .CK(debug_c_c), 
            .Q(count[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i29.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i1 (.D(quadA_delayed_c[0]), .CK(debug_c_c), .Q(quadA_delayed[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i2 (.D(quadA_delayed[1]), .CK(debug_c_c), .Q(quadA_delayed_c[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i2.GSR = "ENABLED";
    CCU2D add_1684_5 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[2]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[3]), .D1(GND_net), .CIN(n26440), .COUT(n26441), 
          .S0(n100[2]), .S1(n100[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_5.INIT0 = 16'h6969;
    defparam add_1684_5.INIT1 = 16'h6969;
    defparam add_1684_5.INJECT1_0 = "NO";
    defparam add_1684_5.INJECT1_1 = "NO";
    LUT4 i2_2_lut (.A(quadB_delayed[2]), .B(quadA_delayed_c[2]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(18[22:95])
    defparam i2_2_lut.init = 16'h6666;
    CCU2D add_1684_3 (.A0(quadA_delayed[1]), .B0(quadB_delayed[2]), .C0(count[0]), 
          .D0(GND_net), .A1(quadA_delayed[1]), .B1(quadB_delayed[2]), 
          .C1(count[1]), .D1(GND_net), .CIN(n26439), .COUT(n26440), 
          .S0(n4358[0]), .S1(n100[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1684_3.INIT0 = 16'h9696;
    defparam add_1684_3.INIT1 = 16'h6969;
    defparam add_1684_3.INJECT1_0 = "NO";
    defparam add_1684_3.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0110000) 
//

module \ArmPeripheral(axis_haddr=8'b0110000)  (read_value, debug_c_c, n2858, 
            n31512, n3922, VCC_net, GND_net, Stepper_A_nFault_c, \read_size[0] , 
            n29258, Stepper_A_M0_c_0, databus, limit_latched, prev_limit_latched, 
            n9331, prev_select, n31445, Stepper_A_M1_c_1, \register_addr[0] , 
            \register_addr[1] , n224, n32, n32_adj_1, prev_step_clk, 
            step_clk, n31419, n22, prev_step_clk_adj_2, n34, step_clk_adj_3, 
            n31421, n24, n31428, \register_addr[5] , n31497, n29271, 
            n31576, n27442, \read_size[2] , n29257, Stepper_A_M2_c_2, 
            Stepper_A_Dir_c, Stepper_A_En_c, \control_reg[7] , n12211, 
            Stepper_A_Step_c, limit_c_3, n8654, n31410, n8402, n8368, 
            n16843) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    input n2858;
    input n31512;
    input [31:0]n3922;
    input VCC_net;
    input GND_net;
    input Stepper_A_nFault_c;
    output \read_size[0] ;
    input n29258;
    output Stepper_A_M0_c_0;
    input [31:0]databus;
    output limit_latched;
    output prev_limit_latched;
    input n9331;
    output prev_select;
    input n31445;
    output Stepper_A_M1_c_1;
    input \register_addr[0] ;
    input \register_addr[1] ;
    output [31:0]n224;
    input n32;
    input n32_adj_1;
    input prev_step_clk;
    input step_clk;
    output n31419;
    output n22;
    input prev_step_clk_adj_2;
    input n34;
    input step_clk_adj_3;
    output n31421;
    output n24;
    input n31428;
    input \register_addr[5] ;
    input n31497;
    input n29271;
    input n31576;
    output n27442;
    output \read_size[2] ;
    input n29257;
    output Stepper_A_M2_c_2;
    output Stepper_A_Dir_c;
    output Stepper_A_En_c;
    output \control_reg[7] ;
    input n12211;
    output Stepper_A_Step_c;
    input limit_c_3;
    input n8654;
    input n31410;
    output n8402;
    output n8368;
    input n16843;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire n49, n41, n60, n54, n42, n62, n52, n38, n58, n50, 
        n56, n46, n9556, n29692, fault_latched, n13943, prev_step_clk_c, 
        step_clk_c, n182;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n29699, n29700;
    wire [31:0]n100;
    
    wire n29731, n29701, n26835, n26834, n31417, n22_c, n26833, 
        n26832, n26831, n26830, n26829, n26828, n26827, n26826, 
        n26825, n26824, n26823, n26822, n26821, n26820, n29729, 
        n29730, n29690, n29691;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire int_step;
    wire [7:0]n8653;
    wire [31:0]n7371;
    
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[0]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52), .C(n38), .D(steps_reg[18]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[7]), .B(steps_reg[9]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[26]), .B(n56), .C(n46), .D(steps_reg[29]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    FD1P3IX read_value__i0 (.D(n29692), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i22_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[25]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[10]), .B(steps_reg[22]), .C(steps_reg[20]), 
         .D(steps_reg[3]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[5]), .B(steps_reg[6]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[28]), .C(steps_reg[13]), 
         .D(steps_reg[30]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[2]), .B(steps_reg[8]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    FD1S3IX steps_reg__i0 (.D(n3922[0]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_A_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n29258), .SP(n2858), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3IX control_reg_i1 (.D(databus[0]), .SP(n13943), .CD(n31512), 
            .CK(debug_c_c), .Q(Stepper_A_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk_c), .CK(debug_c_c), .Q(prev_step_clk_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i0 (.D(databus[0]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n31445), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3922[31]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3922[30]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3922[29]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3922[28]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3922[27]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3922[26]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3922[25]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3922[24]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3922[23]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3922[22]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3922[21]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3922[20]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3922[19]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3922[18]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3922[17]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3922[16]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3922[15]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3922[14]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3922[13]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3922[12]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3922[11]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3922[10]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3922[9]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3922[8]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3922[7]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3922[6]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3922[5]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3922[4]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3922[3]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3922[2]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3922[1]), .CK(debug_c_c), .CD(n31512), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 i22139_3_lut (.A(Stepper_A_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n29699)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22139_3_lut.init = 16'hcaca;
    LUT4 i22140_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n29700)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22140_3_lut.init = 16'hcaca;
    LUT4 i14872_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14872_4_lut.init = 16'hc088;
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    LUT4 i14873_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14873_4_lut.init = 16'hc088;
    LUT4 i14874_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14874_4_lut.init = 16'hc088;
    LUT4 i14875_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14875_4_lut.init = 16'hc088;
    LUT4 i14876_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14876_4_lut.init = 16'hc088;
    LUT4 i14877_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n100[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14877_4_lut.init = 16'hc088;
    LUT4 i14878_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14878_4_lut.init = 16'hc088;
    LUT4 i14879_4_lut (.A(div_factor_reg[24]), .B(\register_addr[1] ), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14879_4_lut.init = 16'hc088;
    LUT4 i14880_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n100[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14880_4_lut.init = 16'hc088;
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n100[26]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n100[23]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n100[20]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n100[7]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n29731), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n29701), .SP(n2858), .CD(n9556), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i14881_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14881_4_lut.init = 16'hc088;
    LUT4 i14882_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14882_4_lut.init = 16'hc088;
    LUT4 i14883_4_lut (.A(div_factor_reg[20]), .B(\register_addr[1] ), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n100[20])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14883_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26835), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26834), .COUT(n26835), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_273 (.A(n32), .B(prev_step_clk_c), .C(step_clk_c), 
         .Z(n31417)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_273.init = 16'h2020;
    LUT4 i14884_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14884_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_4_lut (.A(n32), .B(prev_step_clk_c), .C(step_clk_c), 
         .D(n31512), .Z(n22_c)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut.init = 16'h002c;
    LUT4 i14885_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14885_4_lut.init = 16'hc088;
    LUT4 i14886_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14886_4_lut.init = 16'hc088;
    LUT4 i2_3_lut_rep_275 (.A(n32_adj_1), .B(prev_step_clk), .C(step_clk), 
         .Z(n31419)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_275.init = 16'h2020;
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26833), .COUT(n26834), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut_adj_1 (.A(n32_adj_1), .B(prev_step_clk), .C(step_clk), 
         .D(n31512), .Z(n22)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_1.init = 16'h002c;
    LUT4 i14887_4_lut (.A(div_factor_reg[16]), .B(\register_addr[1] ), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n100[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14887_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26832), .COUT(n26833), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    LUT4 i14888_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14888_4_lut.init = 16'hc088;
    LUT4 i14889_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14889_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26831), .COUT(n26832), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    LUT4 i14890_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14890_4_lut.init = 16'hc088;
    LUT4 i14891_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14891_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26830), .COUT(n26831), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26829), .COUT(n26830), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    LUT4 i14892_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14892_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26828), .COUT(n26829), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26827), .COUT(n26828), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26826), .COUT(n26827), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26825), .COUT(n26826), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_277 (.A(prev_step_clk_adj_2), .B(n34), .C(step_clk_adj_3), 
         .Z(n31421)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_277.init = 16'h4040;
    LUT4 i14893_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14893_4_lut.init = 16'hc088;
    LUT4 i14894_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14894_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26824), .COUT(n26825), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26823), .COUT(n26824), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    LUT4 i14895_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14895_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26822), .COUT(n26823), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut_adj_2 (.A(prev_step_clk_adj_2), .B(n34), .C(step_clk_adj_3), 
         .D(n31512), .Z(n24)) /* synthesis lut_function=(!(A (C+(D))+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_2.init = 16'h004a;
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26821), .COUT(n26822), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26820), .COUT(n26821), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk_c), .D1(prev_step_clk_c), 
          .COUT(n26820), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(n31428), .B(n31512), .C(\register_addr[5] ), .D(n31497), 
         .Z(n9556)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i2_4_lut.init = 16'h0222;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n31445), .B(prev_select), .C(n29271), 
         .D(n31576), .Z(n13943)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n27442)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    PFUMX i22171 (.BLUT(n29729), .ALUT(n29730), .C0(\register_addr[0] ), 
          .Z(n29731));
    FD1P3AX read_size__i2 (.D(n29257), .SP(n2858), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    PFUMX i22132 (.BLUT(n29690), .ALUT(n29691), .C0(\register_addr[1] ), 
          .Z(n29692));
    PFUMX i22141 (.BLUT(n29699), .ALUT(n29700), .C0(\register_addr[1] ), 
          .Z(n29701));
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n13943), .PD(n31512), 
            .CK(debug_c_c), .Q(Stepper_A_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n13943), .CD(n31512), 
            .CK(debug_c_c), .Q(Stepper_A_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n13943), .PD(n31512), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n13943), .CD(n31512), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n13943), .PD(n31512), 
            .CK(debug_c_c), .Q(Stepper_A_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n13943), .PD(n31512), 
            .CK(debug_c_c), .Q(Stepper_A_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n13943), .CD(n12211), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n9331), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n9331), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n9331), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n9331), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n9331), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n9331), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n9331), .PD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n9331), .CD(n31512), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_A_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 i22169_3_lut (.A(Stepper_A_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n29729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22169_3_lut.init = 16'hcaca;
    LUT4 i22170_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n29730)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22170_3_lut.init = 16'hcaca;
    FD1P3AX int_step_182 (.D(n31417), .SP(n22_c), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 i118_1_lut (.A(limit_c_3), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i22130_3_lut (.A(Stepper_A_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n29690)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22130_3_lut.init = 16'hcaca;
    LUT4 i14871_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n8653[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14871_2_lut.init = 16'h2222;
    LUT4 mux_2002_i4_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), .C(\register_addr[0] ), 
         .Z(n7371[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_2002_i4_3_lut.init = 16'hcaca;
    LUT4 i14870_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n8653[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14870_2_lut.init = 16'h2222;
    LUT4 mux_2002_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n7371[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_2002_i5_3_lut.init = 16'hcaca;
    LUT4 i14869_2_lut (.A(Stepper_A_Dir_c), .B(\register_addr[0] ), .Z(n8653[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14869_2_lut.init = 16'h2222;
    LUT4 mux_2002_i6_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), .C(\register_addr[0] ), 
         .Z(n7371[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_2002_i6_3_lut.init = 16'hcaca;
    LUT4 i14868_2_lut (.A(Stepper_A_En_c), .B(\register_addr[0] ), .Z(n8653[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14868_2_lut.init = 16'h2222;
    LUT4 i22131_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n29691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22131_3_lut.init = 16'hcaca;
    LUT4 mux_2002_i7_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n7371[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_2002_i7_3_lut.init = 16'hcaca;
    LUT4 mux_2002_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n7371[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_2002_i8_3_lut.init = 16'hcaca;
    PFUMX mux_2006_i4 (.BLUT(n8653[3]), .ALUT(n7371[3]), .C0(\register_addr[1] ), 
          .Z(n100[3]));
    PFUMX mux_2006_i5 (.BLUT(n8653[4]), .ALUT(n7371[4]), .C0(\register_addr[1] ), 
          .Z(n100[4]));
    PFUMX mux_2006_i6 (.BLUT(n8653[5]), .ALUT(n7371[5]), .C0(\register_addr[1] ), 
          .Z(n100[5]));
    PFUMX mux_2006_i7 (.BLUT(n8653[6]), .ALUT(n7371[6]), .C0(\register_addr[1] ), 
          .Z(n100[6]));
    PFUMX mux_2006_i8 (.BLUT(n8654), .ALUT(n7371[7]), .C0(\register_addr[1] ), 
          .Z(n100[7]));
    ClockDivider_U9 step_clk_gen (.GND_net(GND_net), .step_clk(step_clk_c), 
            .debug_c_c(debug_c_c), .n31512(n31512), .n31410(n31410), .div_factor_reg({div_factor_reg}), 
            .n8402(n8402), .n8368(n8368), .n16843(n16843)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U9
//

module ClockDivider_U9 (GND_net, step_clk, debug_c_c, n31512, n31410, 
            div_factor_reg, n8402, n8368, n16843) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output step_clk;
    input debug_c_c;
    input n31512;
    input n31410;
    input [31:0]div_factor_reg;
    output n8402;
    output n8368;
    input n16843;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n26551;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n26552, n26550, n26549, n26548, n8333, n26547, n26546, 
        n26545, n26544, n26955;
    wire [31:0]n134;
    
    wire n26954, n26953, n26952, n26951, n26543, n26542, n26950, 
        n26949, n26948, n26947, n26946, n26945, n26944, n26943, 
        n26942, n26941, n26940, n27115, n27114, n27113, n27112, 
        n27111, n27110, n27109, n27108, n27107, n27106, n26541, 
        n27105, n26540, n26539;
    wire [31:0]n40;
    
    wire n26538, n26537, n26536, n26535, n27104, n26534, n26533, 
        n27103, n26532, n26531, n26530, n26529, n26528, n26527, 
        n26526, n27102, n26525, n26524, n27101, n27100, n26771, 
        n26770, n26769, n26768, n26767, n26766, n26765, n26764, 
        n26763, n26762, n26761, n26760, n26759, n26758, n26757, 
        n26756, n26555, n26554, n26553;
    
    CCU2D sub_2079_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26551), .COUT(n26552));
    defparam sub_2079_add_2_25.INIT0 = 16'h5999;
    defparam sub_2079_add_2_25.INIT1 = 16'h5999;
    defparam sub_2079_add_2_25.INJECT1_0 = "NO";
    defparam sub_2079_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2079_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26550), .COUT(n26551));
    defparam sub_2079_add_2_23.INIT0 = 16'h5999;
    defparam sub_2079_add_2_23.INIT1 = 16'h5999;
    defparam sub_2079_add_2_23.INJECT1_0 = "NO";
    defparam sub_2079_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2079_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26549), .COUT(n26550));
    defparam sub_2079_add_2_21.INIT0 = 16'h5999;
    defparam sub_2079_add_2_21.INIT1 = 16'h5999;
    defparam sub_2079_add_2_21.INJECT1_0 = "NO";
    defparam sub_2079_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2079_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26548), .COUT(n26549));
    defparam sub_2079_add_2_19.INIT0 = 16'h5999;
    defparam sub_2079_add_2_19.INIT1 = 16'h5999;
    defparam sub_2079_add_2_19.INJECT1_0 = "NO";
    defparam sub_2079_add_2_19.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n8333), .CK(debug_c_c), .CD(n31512), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2079_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26547), .COUT(n26548));
    defparam sub_2079_add_2_17.INIT0 = 16'h5999;
    defparam sub_2079_add_2_17.INIT1 = 16'h5999;
    defparam sub_2079_add_2_17.INJECT1_0 = "NO";
    defparam sub_2079_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2079_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26546), .COUT(n26547));
    defparam sub_2079_add_2_15.INIT0 = 16'h5999;
    defparam sub_2079_add_2_15.INIT1 = 16'h5999;
    defparam sub_2079_add_2_15.INJECT1_0 = "NO";
    defparam sub_2079_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2079_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26545), .COUT(n26546));
    defparam sub_2079_add_2_13.INIT0 = 16'h5999;
    defparam sub_2079_add_2_13.INIT1 = 16'h5999;
    defparam sub_2079_add_2_13.INJECT1_0 = "NO";
    defparam sub_2079_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2079_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26544), .COUT(n26545));
    defparam sub_2079_add_2_11.INIT0 = 16'h5999;
    defparam sub_2079_add_2_11.INIT1 = 16'h5999;
    defparam sub_2079_add_2_11.INJECT1_0 = "NO";
    defparam sub_2079_add_2_11.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26955), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_33.INIT1 = 16'h0000;
    defparam count_2677_add_4_33.INJECT1_0 = "NO";
    defparam count_2677_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26954), .COUT(n26955), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_31.INJECT1_0 = "NO";
    defparam count_2677_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26953), .COUT(n26954), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_29.INJECT1_0 = "NO";
    defparam count_2677_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26952), .COUT(n26953), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_27.INJECT1_0 = "NO";
    defparam count_2677_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26951), .COUT(n26952), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_25.INJECT1_0 = "NO";
    defparam count_2677_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_2079_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26543), .COUT(n26544));
    defparam sub_2079_add_2_9.INIT0 = 16'h5999;
    defparam sub_2079_add_2_9.INIT1 = 16'h5999;
    defparam sub_2079_add_2_9.INJECT1_0 = "NO";
    defparam sub_2079_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2079_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26542), .COUT(n26543));
    defparam sub_2079_add_2_7.INIT0 = 16'h5999;
    defparam sub_2079_add_2_7.INIT1 = 16'h5999;
    defparam sub_2079_add_2_7.INJECT1_0 = "NO";
    defparam sub_2079_add_2_7.INJECT1_1 = "NO";
    FD1S3IX count_2677__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i0.GSR = "ENABLED";
    CCU2D count_2677_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26950), .COUT(n26951), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_23.INJECT1_0 = "NO";
    defparam count_2677_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26949), .COUT(n26950), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_21.INJECT1_0 = "NO";
    defparam count_2677_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26948), .COUT(n26949), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_19.INJECT1_0 = "NO";
    defparam count_2677_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26947), .COUT(n26948), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_17.INJECT1_0 = "NO";
    defparam count_2677_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26946), .COUT(n26947), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_15.INJECT1_0 = "NO";
    defparam count_2677_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26945), .COUT(n26946), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_13.INJECT1_0 = "NO";
    defparam count_2677_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26944), .COUT(n26945), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_11.INJECT1_0 = "NO";
    defparam count_2677_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26943), .COUT(n26944), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_9.INJECT1_0 = "NO";
    defparam count_2677_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26942), .COUT(n26943), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_7.INJECT1_0 = "NO";
    defparam count_2677_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26941), .COUT(n26942), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_5.INJECT1_0 = "NO";
    defparam count_2677_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26940), .COUT(n26941), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2677_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2677_add_4_3.INJECT1_0 = "NO";
    defparam count_2677_add_4_3.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27115), .S1(n8402));
    defparam sub_2082_add_2_33.INIT0 = 16'hf555;
    defparam sub_2082_add_2_33.INIT1 = 16'h0000;
    defparam sub_2082_add_2_33.INJECT1_0 = "NO";
    defparam sub_2082_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27114), .COUT(n27115));
    defparam sub_2082_add_2_31.INIT0 = 16'hf555;
    defparam sub_2082_add_2_31.INIT1 = 16'hf555;
    defparam sub_2082_add_2_31.INJECT1_0 = "NO";
    defparam sub_2082_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27113), .COUT(n27114));
    defparam sub_2082_add_2_29.INIT0 = 16'hf555;
    defparam sub_2082_add_2_29.INIT1 = 16'hf555;
    defparam sub_2082_add_2_29.INJECT1_0 = "NO";
    defparam sub_2082_add_2_29.INJECT1_1 = "NO";
    CCU2D count_2677_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26940), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677_add_4_1.INIT0 = 16'hF000;
    defparam count_2677_add_4_1.INIT1 = 16'h0555;
    defparam count_2677_add_4_1.INJECT1_0 = "NO";
    defparam count_2677_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27112), .COUT(n27113));
    defparam sub_2082_add_2_27.INIT0 = 16'hf555;
    defparam sub_2082_add_2_27.INIT1 = 16'hf555;
    defparam sub_2082_add_2_27.INJECT1_0 = "NO";
    defparam sub_2082_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27111), .COUT(n27112));
    defparam sub_2082_add_2_25.INIT0 = 16'hf555;
    defparam sub_2082_add_2_25.INIT1 = 16'hf555;
    defparam sub_2082_add_2_25.INJECT1_0 = "NO";
    defparam sub_2082_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27110), .COUT(n27111));
    defparam sub_2082_add_2_23.INIT0 = 16'hf555;
    defparam sub_2082_add_2_23.INIT1 = 16'hf555;
    defparam sub_2082_add_2_23.INJECT1_0 = "NO";
    defparam sub_2082_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27109), .COUT(n27110));
    defparam sub_2082_add_2_21.INIT0 = 16'hf555;
    defparam sub_2082_add_2_21.INIT1 = 16'hf555;
    defparam sub_2082_add_2_21.INJECT1_0 = "NO";
    defparam sub_2082_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27108), .COUT(n27109));
    defparam sub_2082_add_2_19.INIT0 = 16'hf555;
    defparam sub_2082_add_2_19.INIT1 = 16'hf555;
    defparam sub_2082_add_2_19.INJECT1_0 = "NO";
    defparam sub_2082_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27107), .COUT(n27108));
    defparam sub_2082_add_2_17.INIT0 = 16'hf555;
    defparam sub_2082_add_2_17.INIT1 = 16'hf555;
    defparam sub_2082_add_2_17.INJECT1_0 = "NO";
    defparam sub_2082_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27106), .COUT(n27107));
    defparam sub_2082_add_2_15.INIT0 = 16'hf555;
    defparam sub_2082_add_2_15.INIT1 = 16'hf555;
    defparam sub_2082_add_2_15.INJECT1_0 = "NO";
    defparam sub_2082_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2079_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26541), .COUT(n26542));
    defparam sub_2079_add_2_5.INIT0 = 16'h5999;
    defparam sub_2079_add_2_5.INIT1 = 16'h5999;
    defparam sub_2079_add_2_5.INJECT1_0 = "NO";
    defparam sub_2079_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27105), .COUT(n27106));
    defparam sub_2082_add_2_13.INIT0 = 16'hf555;
    defparam sub_2082_add_2_13.INIT1 = 16'hf555;
    defparam sub_2082_add_2_13.INJECT1_0 = "NO";
    defparam sub_2082_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2079_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26540), .COUT(n26541));
    defparam sub_2079_add_2_3.INIT0 = 16'h5999;
    defparam sub_2079_add_2_3.INIT1 = 16'h5999;
    defparam sub_2079_add_2_3.INJECT1_0 = "NO";
    defparam sub_2079_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2079_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n26540));
    defparam sub_2079_add_2_1.INIT0 = 16'h0000;
    defparam sub_2079_add_2_1.INIT1 = 16'h5999;
    defparam sub_2079_add_2_1.INJECT1_0 = "NO";
    defparam sub_2079_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26539), .S1(n8368));
    defparam sub_2081_add_2_33.INIT0 = 16'h5999;
    defparam sub_2081_add_2_33.INIT1 = 16'h0000;
    defparam sub_2081_add_2_33.INJECT1_0 = "NO";
    defparam sub_2081_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26538), .COUT(n26539));
    defparam sub_2081_add_2_31.INIT0 = 16'h5999;
    defparam sub_2081_add_2_31.INIT1 = 16'h5999;
    defparam sub_2081_add_2_31.INJECT1_0 = "NO";
    defparam sub_2081_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26537), .COUT(n26538));
    defparam sub_2081_add_2_29.INIT0 = 16'h5999;
    defparam sub_2081_add_2_29.INIT1 = 16'h5999;
    defparam sub_2081_add_2_29.INJECT1_0 = "NO";
    defparam sub_2081_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26536), .COUT(n26537));
    defparam sub_2081_add_2_27.INIT0 = 16'h5999;
    defparam sub_2081_add_2_27.INIT1 = 16'h5999;
    defparam sub_2081_add_2_27.INJECT1_0 = "NO";
    defparam sub_2081_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26535), .COUT(n26536));
    defparam sub_2081_add_2_25.INIT0 = 16'h5999;
    defparam sub_2081_add_2_25.INIT1 = 16'h5999;
    defparam sub_2081_add_2_25.INJECT1_0 = "NO";
    defparam sub_2081_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27104), .COUT(n27105));
    defparam sub_2082_add_2_11.INIT0 = 16'hf555;
    defparam sub_2082_add_2_11.INIT1 = 16'hf555;
    defparam sub_2082_add_2_11.INJECT1_0 = "NO";
    defparam sub_2082_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26534), .COUT(n26535));
    defparam sub_2081_add_2_23.INIT0 = 16'h5999;
    defparam sub_2081_add_2_23.INIT1 = 16'h5999;
    defparam sub_2081_add_2_23.INJECT1_0 = "NO";
    defparam sub_2081_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26533), .COUT(n26534));
    defparam sub_2081_add_2_21.INIT0 = 16'h5999;
    defparam sub_2081_add_2_21.INIT1 = 16'h5999;
    defparam sub_2081_add_2_21.INJECT1_0 = "NO";
    defparam sub_2081_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27103), .COUT(n27104));
    defparam sub_2082_add_2_9.INIT0 = 16'hf555;
    defparam sub_2082_add_2_9.INIT1 = 16'hf555;
    defparam sub_2082_add_2_9.INJECT1_0 = "NO";
    defparam sub_2082_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26532), .COUT(n26533));
    defparam sub_2081_add_2_19.INIT0 = 16'h5999;
    defparam sub_2081_add_2_19.INIT1 = 16'h5999;
    defparam sub_2081_add_2_19.INJECT1_0 = "NO";
    defparam sub_2081_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26531), .COUT(n26532));
    defparam sub_2081_add_2_17.INIT0 = 16'h5999;
    defparam sub_2081_add_2_17.INIT1 = 16'h5999;
    defparam sub_2081_add_2_17.INJECT1_0 = "NO";
    defparam sub_2081_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26530), .COUT(n26531));
    defparam sub_2081_add_2_15.INIT0 = 16'h5999;
    defparam sub_2081_add_2_15.INIT1 = 16'h5999;
    defparam sub_2081_add_2_15.INJECT1_0 = "NO";
    defparam sub_2081_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26529), .COUT(n26530));
    defparam sub_2081_add_2_13.INIT0 = 16'h5999;
    defparam sub_2081_add_2_13.INIT1 = 16'h5999;
    defparam sub_2081_add_2_13.INJECT1_0 = "NO";
    defparam sub_2081_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26528), .COUT(n26529));
    defparam sub_2081_add_2_11.INIT0 = 16'h5999;
    defparam sub_2081_add_2_11.INIT1 = 16'h5999;
    defparam sub_2081_add_2_11.INJECT1_0 = "NO";
    defparam sub_2081_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26527), .COUT(n26528));
    defparam sub_2081_add_2_9.INIT0 = 16'h5999;
    defparam sub_2081_add_2_9.INIT1 = 16'h5999;
    defparam sub_2081_add_2_9.INJECT1_0 = "NO";
    defparam sub_2081_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26526), .COUT(n26527));
    defparam sub_2081_add_2_7.INIT0 = 16'h5999;
    defparam sub_2081_add_2_7.INIT1 = 16'h5999;
    defparam sub_2081_add_2_7.INJECT1_0 = "NO";
    defparam sub_2081_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27102), .COUT(n27103));
    defparam sub_2082_add_2_7.INIT0 = 16'hf555;
    defparam sub_2082_add_2_7.INIT1 = 16'hf555;
    defparam sub_2082_add_2_7.INJECT1_0 = "NO";
    defparam sub_2082_add_2_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_2081_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26525), .COUT(n26526));
    defparam sub_2081_add_2_5.INIT0 = 16'h5999;
    defparam sub_2081_add_2_5.INIT1 = 16'h5999;
    defparam sub_2081_add_2_5.INJECT1_0 = "NO";
    defparam sub_2081_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n26524), .COUT(n26525));
    defparam sub_2081_add_2_3.INIT0 = 16'h5999;
    defparam sub_2081_add_2_3.INIT1 = 16'h5999;
    defparam sub_2081_add_2_3.INJECT1_0 = "NO";
    defparam sub_2081_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2081_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n26524));
    defparam sub_2081_add_2_1.INIT0 = 16'h0000;
    defparam sub_2081_add_2_1.INIT1 = 16'h5999;
    defparam sub_2081_add_2_1.INJECT1_0 = "NO";
    defparam sub_2081_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27101), .COUT(n27102));
    defparam sub_2082_add_2_5.INIT0 = 16'hf555;
    defparam sub_2082_add_2_5.INIT1 = 16'hf555;
    defparam sub_2082_add_2_5.INJECT1_0 = "NO";
    defparam sub_2082_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27100), .COUT(n27101));
    defparam sub_2082_add_2_3.INIT0 = 16'hf555;
    defparam sub_2082_add_2_3.INIT1 = 16'hf555;
    defparam sub_2082_add_2_3.INJECT1_0 = "NO";
    defparam sub_2082_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2082_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27100));
    defparam sub_2082_add_2_1.INIT0 = 16'h0000;
    defparam sub_2082_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2082_add_2_1.INJECT1_0 = "NO";
    defparam sub_2082_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n31410), .CD(n16843), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n31410), .PD(n16843), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26771), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26770), .COUT(n26771), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26769), .COUT(n26770), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26768), .COUT(n26769), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26767), .COUT(n26768), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26766), .COUT(n26767), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26765), .COUT(n26766), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26764), .COUT(n26765), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26763), .COUT(n26764), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26762), .COUT(n26763), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26761), .COUT(n26762), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26760), .COUT(n26761), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26759), .COUT(n26760), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26758), .COUT(n26759), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26757), .COUT(n26758), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n26756), .COUT(n26757), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n26756), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    FD1S3IX count_2677__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i1.GSR = "ENABLED";
    FD1S3IX count_2677__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i2.GSR = "ENABLED";
    FD1S3IX count_2677__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i3.GSR = "ENABLED";
    FD1S3IX count_2677__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i4.GSR = "ENABLED";
    FD1S3IX count_2677__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i5.GSR = "ENABLED";
    FD1S3IX count_2677__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i6.GSR = "ENABLED";
    FD1S3IX count_2677__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i7.GSR = "ENABLED";
    FD1S3IX count_2677__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i8.GSR = "ENABLED";
    FD1S3IX count_2677__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i9.GSR = "ENABLED";
    FD1S3IX count_2677__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i10.GSR = "ENABLED";
    FD1S3IX count_2677__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i11.GSR = "ENABLED";
    FD1S3IX count_2677__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i12.GSR = "ENABLED";
    FD1S3IX count_2677__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i13.GSR = "ENABLED";
    FD1S3IX count_2677__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i14.GSR = "ENABLED";
    FD1S3IX count_2677__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i15.GSR = "ENABLED";
    FD1S3IX count_2677__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i16.GSR = "ENABLED";
    FD1S3IX count_2677__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i17.GSR = "ENABLED";
    FD1S3IX count_2677__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i18.GSR = "ENABLED";
    FD1S3IX count_2677__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i19.GSR = "ENABLED";
    FD1S3IX count_2677__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i20.GSR = "ENABLED";
    FD1S3IX count_2677__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i21.GSR = "ENABLED";
    FD1S3IX count_2677__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i22.GSR = "ENABLED";
    FD1S3IX count_2677__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i23.GSR = "ENABLED";
    FD1S3IX count_2677__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i24.GSR = "ENABLED";
    FD1S3IX count_2677__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i25.GSR = "ENABLED";
    FD1S3IX count_2677__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i26.GSR = "ENABLED";
    FD1S3IX count_2677__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i27.GSR = "ENABLED";
    FD1S3IX count_2677__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i28.GSR = "ENABLED";
    FD1S3IX count_2677__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i29.GSR = "ENABLED";
    FD1S3IX count_2677__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i30.GSR = "ENABLED";
    FD1S3IX count_2677__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n31410), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2677__i31.GSR = "ENABLED";
    CCU2D sub_2079_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n26555), .S1(n8333));
    defparam sub_2079_add_2_33.INIT0 = 16'h5555;
    defparam sub_2079_add_2_33.INIT1 = 16'h0000;
    defparam sub_2079_add_2_33.INJECT1_0 = "NO";
    defparam sub_2079_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2079_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26554), .COUT(n26555));
    defparam sub_2079_add_2_31.INIT0 = 16'h5999;
    defparam sub_2079_add_2_31.INIT1 = 16'h5999;
    defparam sub_2079_add_2_31.INJECT1_0 = "NO";
    defparam sub_2079_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2079_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26553), .COUT(n26554));
    defparam sub_2079_add_2_29.INIT0 = 16'h5999;
    defparam sub_2079_add_2_29.INIT1 = 16'h5999;
    defparam sub_2079_add_2_29.INJECT1_0 = "NO";
    defparam sub_2079_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2079_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n26552), .COUT(n26553));
    defparam sub_2079_add_2_27.INIT0 = 16'h5999;
    defparam sub_2079_add_2_27.INIT1 = 16'h5999;
    defparam sub_2079_add_2_27.INJECT1_0 = "NO";
    defparam sub_2079_add_2_27.INJECT1_1 = "NO";
    
endmodule

// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.4.1.213
// Netlist written on Sat May 14 07:35:11 2016
//
// Verilog Description of module UniboardTop
//

module UniboardTop (uart_rx, uart_tx, status_led, clk_12MHz, Stepper_X_Step, 
            Stepper_X_Dir, Stepper_X_M0, Stepper_X_M1, Stepper_X_M2, 
            Stepper_X_En, Stepper_X_nFault, Stepper_Y_Step, Stepper_Y_Dir, 
            Stepper_Y_M0, Stepper_Y_M1, Stepper_Y_M2, Stepper_Y_En, 
            Stepper_Y_nFault, Stepper_Z_Step, Stepper_Z_Dir, Stepper_Z_M0, 
            Stepper_Z_M1, Stepper_Z_M2, Stepper_Z_En, Stepper_Z_nFault, 
            Stepper_A_Step, Stepper_A_Dir, Stepper_A_M0, Stepper_A_M1, 
            Stepper_A_M2, Stepper_A_En, Stepper_A_nFault, limit, expansion1, 
            expansion2, expansion3, expansion4, expansion5, signal_light, 
            encoder_ra, encoder_rb, encoder_ri, encoder_la, encoder_lb, 
            encoder_li, rc_ch1, rc_ch2, rc_ch3, rc_ch4, rc_ch7, 
            rc_ch8, motor_pwm_l, motor_pwm_r, xbee_pause, debug) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(362[8:19])
    input uart_rx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[13:20])
    output uart_tx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[14:21])
    output [2:0]status_led;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    input clk_12MHz;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    output Stepper_X_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(368[17:31])
    output Stepper_X_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:30])
    output Stepper_X_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:29])
    output Stepper_X_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    output Stepper_X_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    output Stepper_X_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    input Stepper_X_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[16:32])
    output Stepper_Y_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(376[17:31])
    output Stepper_Y_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:30])
    output Stepper_Y_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:29])
    output Stepper_Y_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    output Stepper_Y_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    output Stepper_Y_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    input Stepper_Y_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[16:32])
    output Stepper_Z_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(384[17:31])
    output Stepper_Z_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:30])
    output Stepper_Z_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:29])
    output Stepper_Z_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    output Stepper_Z_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    output Stepper_Z_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    input Stepper_Z_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[16:32])
    output Stepper_A_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(392[17:31])
    output Stepper_A_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:30])
    output Stepper_A_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:29])
    output Stepper_A_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    output Stepper_A_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    output Stepper_A_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    input Stepper_A_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[16:32])
    input [3:0]limit;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    output expansion1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[14:24])
    output expansion2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    output expansion3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    inout expansion4;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[13:23])
    input expansion5 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    output signal_light;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[14:26])
    input encoder_ra;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(408[13:23])
    input encoder_rb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    input encoder_ri;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    input encoder_la;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    input encoder_lb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    input encoder_li;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    input rc_ch1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(415[13:19])
    input rc_ch2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    input rc_ch3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    input rc_ch4;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    input rc_ch7;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    input rc_ch8;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    output motor_pwm_l;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(422[14:25])
    output motor_pwm_r;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    input xbee_pause;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[13:23])
    output [8:0]debug;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [127:0]select /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(455[15:21])
    wire [15:0]battery_voltage;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(18[20:35])
    
    wire VCC_net, uart_rx_c, uart_tx_c, Stepper_X_Step_c, Stepper_X_Dir_c, 
        Stepper_X_M0_c_0, Stepper_X_M1_c_1, Stepper_X_M2_c_2, Stepper_X_En_c, 
        Stepper_X_nFault_c, Stepper_Y_Step_c, Stepper_Y_Dir_c, Stepper_Y_M0_c_0, 
        Stepper_Y_M1_c_1, Stepper_Y_M2_c_2, Stepper_Y_En_c, Stepper_Y_nFault_c, 
        Stepper_Z_Step_c, Stepper_Z_Dir_c, Stepper_Z_M0_c_0, Stepper_Z_M1_c_1, 
        Stepper_Z_M2_c_2, Stepper_Z_En_c, Stepper_Z_nFault_c, Stepper_A_Step_c, 
        Stepper_A_Dir_c, Stepper_A_M0_c_0, Stepper_A_M1_c_1, Stepper_A_M2_c_2, 
        Stepper_A_En_c, Stepper_A_nFault_c, limit_c_3, limit_c_2, limit_c_1, 
        limit_c_0, expansion1_c_9, expansion2_c_10, expansion3_c_11, 
        expansion5_c, signal_light_c, encoder_ra_c, encoder_rb_c, encoder_ri_c, 
        encoder_la_c, encoder_lb_c, encoder_li_c, rc_ch1_c, rc_ch2_c, 
        rc_ch3_c, rc_ch4_c, rc_ch7_c, rc_ch8_c, n11013, xbee_pause_c, 
        debug_c_7, debug_c_5, debug_c_4, debug_c_3, debug_c_2, debug_c_0;
    wire [31:0]databus;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(451[14:21])
    wire [2:0]reg_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(452[13:21])
    wire [7:0]register_addr;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    
    wire rw, n30465;
    wire [15:0]reset_count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(458[13:24])
    
    wire timeout_pause;
    wire [31:0]timeout_count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[13:26])
    
    wire prev_uart_rx, n32166, n28061, n13412, n21442, n13, n21445, 
        n14, n21447, n21453, n21455, n13977, n13976, n13975, n13974, 
        n14114, n12, n8, n32135, n8_adj_568, n16516, n16515, n32165, 
        n28053, n32164, n32163, n22;
    wire [7:0]n8575;
    
    wire n44, n32162;
    wire [31:0]n658;
    
    wire n32, n32161, n2, n2_adj_569;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    wire [31:0]databus_out;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(55[13:24])
    
    wire n8_adj_570, n22_adj_571, n14555, n13899, n32_adj_572, n28062, 
        n13885, n8_adj_573, n13118, n32_adj_574;
    wire [31:0]n1414;
    
    wire n24, n5774, n14493, n29948, n44_adj_575, n30470, n8447, 
        n9309, n13769, n21171, n13_adj_576, n21174, n14_adj_577, 
        n21176, n21182, n21184, n8_adj_578, n2_adj_579, n2_adj_580, 
        n12_adj_581, n34, n8_adj_582, n32160, n112, n2_adj_583, 
        n32159, n2_adj_584, n9478;
    wire [31:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(31[13:23])
    wire [2:0]read_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(32[12:21])
    
    wire prev_select, n46, n29194, n8_adj_585, n5, n2_adj_586;
    wire [7:0]\register[0]_adj_959 ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    wire [7:0]read_value_adj_960;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(92[12:22])
    wire [2:0]read_size_adj_961;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(93[12:21])
    
    wire prev_select_adj_596, n64, n27397, n27396, n4;
    wire [15:0]n281;
    
    wire n30019, n29750, n32134, n27395, n29712;
    wire [31:0]n99_adj_1349;
    
    wire n30320, n27394, n27393, n27392, n2_adj_597, n2_adj_598, 
        n14419, n27391, n5_adj_599, n241;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire step_clk, prev_step_clk;
    wire [31:0]read_value_adj_967;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_968;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_634, n52, n4034, n2776, n29920, n302, n30001, 
        n21718, n29947, n32158, n13605, n28140, n28330;
    wire [7:0]n571;
    
    wire n32129, n28333, n13598, n2_adj_635, n8_adj_636, n2_adj_637;
    wire [7:0]control_reg_adj_976;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire step_clk_adj_639, prev_step_clk_adj_640;
    wire [31:0]read_value_adj_979;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_980;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_675, n13588, n52_adj_676, n2_adj_677, n13576, 
        n8_adj_678, n13567, n8_adj_679, n8_adj_680, n2_adj_681, n8_adj_682, 
        n17, n13560, n16, n28331, n15, n13545;
    wire [31:0]n580_adj_998;
    
    wire n8_adj_683, n8_adj_684, n32140, n2769;
    wire [7:0]control_reg_adj_1014;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]div_factor_reg_adj_1015;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg_adj_1016;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire int_step, step_clk_adj_686, prev_step_clk_adj_687;
    wire [31:0]read_value_adj_1017;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_1018;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_722;
    wire [31:0]n224_adj_1021;
    
    wire n2_adj_724, n2_adj_725;
    wire [31:0]n3948;
    
    wire n32138, n13511, n14355, n44_adj_726, n29759, n30260;
    wire [31:0]n580_adj_1036;
    
    wire n8_adj_727, n32157;
    wire [7:0]control_reg_adj_1052;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]div_factor_reg_adj_1053;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg_adj_1054;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire int_step_adj_738;
    wire [31:0]read_value_adj_1055;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_1056;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_773, n19559, n28133;
    wire [31:0]n224_adj_1059;
    
    wire n2_adj_806, n28365, n2_adj_807, n3, n13476;
    wire [31:0]n3862;
    
    wire n2_adj_808, n9, n28141, n28328, n2_adj_809, n30566, qreset;
    wire [31:0]read_value_adj_1092;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(65[13:23])
    wire [2:0]read_size_adj_1093;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(66[12:21])
    
    wire prev_select_adj_844, n41, n29954, n2_adj_845, n8_adj_846;
    wire [31:0]read_value_adj_1100;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(65[13:23])
    wire [2:0]read_size_adj_1101;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(66[12:21])
    
    wire prev_select_adj_881, n178, n3_adj_882, n2_adj_883, n2760;
    wire [7:0]read_value_adj_1116;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(26[12:22])
    wire [2:0]read_size_adj_1117;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(27[12:21])
    
    wire prev_select_adj_893, n18, n6, n14_adj_894, n176, n13_adj_895, 
        n32155, n8_adj_896, n2_adj_897, n30, n29860, n22529, n16718, 
        n30075, n14812, n29544, n30472, n28231, n28144, n42, n40, 
        n38, n1, n29758, n36, n32154, n34_adj_898, n28329, n30_adj_899, 
        n3_adj_900, n29, n26, n32153, n2_adj_901, n8_adj_902, n2_adj_903, 
        n2_adj_904, n29953, n29977, n2_adj_905, n3_adj_906, n8_adj_907, 
        n32152;
    wire [2:0]quadA_delayed_adj_1199;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    wire [2:0]quadB_delayed_adj_1200;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    
    wire n9496, n9485, n9482, n28017, n142, n14271;
    wire [15:0]count_adj_1215;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n27737, n27736;
    wire [15:0]count_adj_1228;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n5_adj_912, n27735, n27734, n27733, n27732, n7822, n27731, 
        n27730, n27729, n27728, n27727, n205;
    wire [15:0]count_adj_1267;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n5_adj_917, n8_adj_918, n7787, n32317, n32316, n32315, 
        n32314, n30546, n30330, n32308, n32306, n30324, n32305, 
        n34068, n30308, n34065, n11961, n30304, n30020, n107;
    wire [3:0]state_adj_1287;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n30302, n32302, n32301, n30270, n2_adj_919, n21617, n32296, 
        n32294, n32293, n32290, n32137, n29883;
    wire [7:0]n8584;
    
    wire n32285, n32284, n32283;
    wire [31:0]n7033;
    
    wire n32282, n32279, n32278, n34066, n30613, n32274, n28222, 
        n34071;
    wire [7:0]n8593;
    
    wire n32267, n32264, n32261, n32258, n32257, n32256;
    wire [31:0]n7347;
    
    wire n32141, n27046, n32253, n32252, n27045, n32251, n5_adj_920, 
        n8_adj_921, n27044, n32245, n27043, n27042, n27041, n8_adj_922, 
        n9_adj_923, n34070, n27040, n27039, n27038, n30463, n27037, 
        n34067, n32235, n32234, n3_adj_924, n2_adj_925, n32233, 
        n32232, n27036, n32231, n3_adj_926, n2_adj_927, n10, n34069, 
        n3_adj_928, n2_adj_929, n10_adj_930, n32227, n34064, n3_adj_931, 
        n32221, n27035, n27034, n32218, n32216, n32215, n32213, 
        n10948, n30615, n30617, n30619, n30621, n32149, n28233, 
        n30623, n28232, n28234, n10947;
    wire [14:0]n66_adj_1469;
    
    wire n27033, n32205, n32204, n32203, n32202, n29983, n32200, 
        n27032, n32199, n32127, n32189, n32187, n8_adj_932, n27031, 
        n32185, n2_adj_933, n8_adj_934, n32182, n28426, n28302, 
        n32181, n32178, n28129, n28132, n32147, n32146, n32145, 
        n32144, n32142, n32172, n29713, n32125, n28407, n12746, 
        n30482, n30474, n32168, n28049, expansion4_out;
    
    VHI i2 (.Z(VCC_net));
    ExpansionGPIO gpio (.read_value({read_value_adj_1116}), .debug_c_c(debug_c_c), 
            .n32162(n32162), .n13598(n13598), .n34066(n34066), .\databus[0] (databus[0]), 
            .\read_size[0] (read_size_adj_1117[0]), .n22529(n22529), .prev_select(prev_select_adj_893), 
            .\select[5] (select[5]), .n10948(n10948), .n10947(n10947), 
            .expansion1_c_9(expansion1_c_9), .n14812(n14812), .expansion2_c_10(expansion2_c_10), 
            .expansion3_c_11(expansion3_c_11), .expansion5_c(expansion5_c), 
            .n32187(n32187), .n32204(n32204), .\register_addr[0] (register_addr[0]), 
            .expansion4_out(expansion4_out), .n32315(n32315), .n32279(n32279), 
            .n32235(n32235), .n302(n302), .n32158(n32158), .rw(rw), 
            .n32172(n32172), .\register_addr[1] (register_addr[1]), .n32282(n32282), 
            .n21617(n21617), .n32278(n32278), .n32146(n32146), .n32147(n32147), 
            .n32306(n32306), .n32216(n32216), .\databus[1] (databus[1]), 
            .\databus[2] (databus[2]), .\databus[3] (databus[3]), .\databus[4] (databus[4]), 
            .\databus[5] (databus[5]), .\databus[6] (databus[6]), .\databus[7] (databus[7]), 
            .n11961(n11961), .n16718(n16718), .n32232(n32232), .\register_addr[3] (register_addr[3]), 
            .n29920(n29920), .\register_addr[2] (register_addr[2]), .n176(n176), 
            .n32185(n32185), .n112(n112), .n28365(n28365)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(694[18] 705[38])
    IFS1P3DX prev_uart_rx_58 (.D(uart_rx_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(battery_voltage[15]), .Q(prev_uart_rx));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam prev_uart_rx_58.GSR = "ENABLED";
    FD1S3AX timeout_pause_60 (.D(n28407), .CK(debug_c_c), .Q(timeout_pause));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_pause_60.GSR = "ENABLED";
    FD1P3AX timeout_count__i0 (.D(n99_adj_1349[0]), .SP(n14355), .CK(debug_c_c), 
            .Q(timeout_count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i0.GSR = "ENABLED";
    CCU2D add_31_9 (.A0(timeout_count[7]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[8]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27034), 
          .COUT(n27035), .S0(n658[7]), .S1(n658[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_9.INIT0 = 16'h5aaa;
    defparam add_31_9.INIT1 = 16'h5aaa;
    defparam add_31_9.INJECT1_0 = "NO";
    defparam add_31_9.INJECT1_1 = "NO";
    CCU2D add_31_7 (.A0(timeout_count[5]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[6]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27033), 
          .COUT(n27034), .S0(n658[5]), .S1(n658[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_7.INIT0 = 16'h5aaa;
    defparam add_31_7.INIT1 = 16'h5aaa;
    defparam add_31_7.INJECT1_0 = "NO";
    defparam add_31_7.INJECT1_1 = "NO";
    LUT4 i2646_1_lut (.A(n7787), .Z(n9309)) /* synthesis lut_function=(!(A)) */ ;
    defparam i2646_1_lut.init = 16'h5555;
    CCU2D reset_count_2657_2658_add_4_9 (.A0(reset_count[7]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[8]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27394), .COUT(n27395), .S0(n66_adj_1469[7]), .S1(n66_adj_1469[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658_add_4_9.INIT0 = 16'hfaaa;
    defparam reset_count_2657_2658_add_4_9.INIT1 = 16'hfaaa;
    defparam reset_count_2657_2658_add_4_9.INJECT1_0 = "NO";
    defparam reset_count_2657_2658_add_4_9.INJECT1_1 = "NO";
    CCU2D reset_count_2657_2658_add_4_7 (.A0(reset_count[5]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[6]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27393), .COUT(n27394), .S0(n66_adj_1469[5]), .S1(n66_adj_1469[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658_add_4_7.INIT0 = 16'hfaaa;
    defparam reset_count_2657_2658_add_4_7.INIT1 = 16'hfaaa;
    defparam reset_count_2657_2658_add_4_7.INJECT1_0 = "NO";
    defparam reset_count_2657_2658_add_4_7.INJECT1_1 = "NO";
    CCU2D reset_count_2657_2658_add_4_5 (.A0(reset_count[3]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[4]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27392), .COUT(n27393), .S0(n66_adj_1469[3]), .S1(n66_adj_1469[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658_add_4_5.INIT0 = 16'hfaaa;
    defparam reset_count_2657_2658_add_4_5.INIT1 = 16'hfaaa;
    defparam reset_count_2657_2658_add_4_5.INJECT1_0 = "NO";
    defparam reset_count_2657_2658_add_4_5.INJECT1_1 = "NO";
    CCU2D reset_count_2657_2658_add_4_3 (.A0(reset_count[1]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[2]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27391), .COUT(n27392), .S0(n66_adj_1469[1]), .S1(n66_adj_1469[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658_add_4_3.INIT0 = 16'hfaaa;
    defparam reset_count_2657_2658_add_4_3.INIT1 = 16'hfaaa;
    defparam reset_count_2657_2658_add_4_3.INJECT1_0 = "NO";
    defparam reset_count_2657_2658_add_4_3.INJECT1_1 = "NO";
    CCU2D reset_count_2657_2658_add_4_1 (.A0(battery_voltage[15]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[0]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .COUT(n27391), .S1(n66_adj_1469[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658_add_4_1.INIT0 = 16'hF000;
    defparam reset_count_2657_2658_add_4_1.INIT1 = 16'h0555;
    defparam reset_count_2657_2658_add_4_1.INJECT1_0 = "NO";
    defparam reset_count_2657_2658_add_4_1.INJECT1_1 = "NO";
    CCU2D add_31_5 (.A0(timeout_count[3]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[4]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27032), 
          .COUT(n27033), .S0(n658[3]), .S1(n658[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_5.INIT0 = 16'h5aaa;
    defparam add_31_5.INIT1 = 16'h5aaa;
    defparam add_31_5.INJECT1_0 = "NO";
    defparam add_31_5.INJECT1_1 = "NO";
    CCU2D add_31_3 (.A0(timeout_count[1]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[2]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27031), 
          .COUT(n27032), .S0(n658[1]), .S1(n658[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_3.INIT0 = 16'h5aaa;
    defparam add_31_3.INIT1 = 16'h5aaa;
    defparam add_31_3.INJECT1_0 = "NO";
    defparam add_31_3.INJECT1_1 = "NO";
    LUT4 Select_4281_i2_2_lut_3_lut_4_lut (.A(n32261), .B(n32168), .C(read_value_adj_1055[5]), 
         .D(rw), .Z(n2_adj_905)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4281_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4282_i2_2_lut_3_lut_4_lut (.A(n32261), .B(n32168), .C(read_value_adj_1055[4]), 
         .D(rw), .Z(n2_adj_883)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4282_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i186_4_lut (.A(n142), .B(reset_count[5]), .C(reset_count[6]), 
         .D(reset_count[4]), .Z(n205)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(458[13:24])
    defparam i186_4_lut.init = 16'hfaea;
    LUT4 Select_4279_i2_2_lut_3_lut_4_lut (.A(n32261), .B(n32168), .C(read_value_adj_1055[7]), 
         .D(rw), .Z(n2_adj_807)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4279_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    CCU2D add_31_1 (.A0(battery_voltage[15]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[0]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .COUT(n27031), .S1(n658[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_1.INIT0 = 16'hF000;
    defparam add_31_1.INIT1 = 16'h5555;
    defparam add_31_1.INJECT1_0 = "NO";
    defparam add_31_1.INJECT1_1 = "NO";
    LUT4 i23032_2_lut (.A(int_step_adj_738), .B(control_reg_adj_1052[3]), 
         .Z(Stepper_A_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i23032_2_lut.init = 16'h9999;
    LUT4 i23030_2_lut (.A(int_step), .B(control_reg_adj_1014[3]), .Z(Stepper_Z_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i23030_2_lut.init = 16'h9999;
    LUT4 Select_4286_i2_2_lut_3_lut_4_lut (.A(n32261), .B(n32168), .C(read_value_adj_1055[0]), 
         .D(rw), .Z(n2_adj_927)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4286_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    IB xbee_pause_pad (.I(xbee_pause), .O(xbee_pause_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[13:23])
    IB rc_ch8_pad (.I(rc_ch8), .O(rc_ch8_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    IB rc_ch7_pad (.I(rc_ch7), .O(rc_ch7_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    IB rc_ch4_pad (.I(rc_ch4), .O(rc_ch4_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    IB rc_ch3_pad (.I(rc_ch3), .O(rc_ch3_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    IB rc_ch2_pad (.I(rc_ch2), .O(rc_ch2_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    IB rc_ch1_pad (.I(rc_ch1), .O(rc_ch1_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(415[13:19])
    IB encoder_li_pad (.I(encoder_li), .O(encoder_li_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    IB encoder_lb_pad (.I(encoder_lb), .O(encoder_lb_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    IB encoder_la_pad (.I(encoder_la), .O(encoder_la_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    IB encoder_ri_pad (.I(encoder_ri), .O(encoder_ri_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    IB encoder_rb_pad (.I(encoder_rb), .O(encoder_rb_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    IB encoder_ra_pad (.I(encoder_ra), .O(encoder_ra_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(408[13:23])
    IB expansion5_pad (.I(expansion5), .O(expansion5_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    IB limit_pad_0 (.I(limit[0]), .O(limit_c_0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB limit_pad_1 (.I(limit[1]), .O(limit_c_1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB limit_pad_2 (.I(limit[2]), .O(limit_c_2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB limit_pad_3 (.I(limit[3]), .O(limit_c_3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(400[19:24])
    IB Stepper_A_nFault_pad (.I(Stepper_A_nFault), .O(Stepper_A_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[16:32])
    IB Stepper_Z_nFault_pad (.I(Stepper_Z_nFault), .O(Stepper_Z_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[16:32])
    IB Stepper_Y_nFault_pad (.I(Stepper_Y_nFault), .O(Stepper_Y_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[16:32])
    IB Stepper_X_nFault_pad (.I(Stepper_X_nFault), .O(Stepper_X_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[16:32])
    IB debug_c_pad (.I(clk_12MHz), .O(debug_c_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    IB uart_rx_pad (.I(uart_rx), .O(uart_rx_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[13:20])
    OB debug_pad_0 (.I(debug_c_0), .O(debug[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_1 (.I(n11013), .O(debug[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_2 (.I(debug_c_2), .O(debug[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_3 (.I(debug_c_3), .O(debug[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_4 (.I(debug_c_4), .O(debug[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_5 (.I(debug_c_5), .O(debug[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_6 (.I(n34065), .O(debug[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_7 (.I(debug_c_7), .O(debug[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB debug_pad_8 (.I(debug_c_c), .O(debug[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(426[19:24])
    OB motor_pwm_r_pad (.I(n11013), .O(motor_pwm_r));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    OB motor_pwm_l_pad (.I(n11013), .O(motor_pwm_l));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(422[14:25])
    OB signal_light_pad (.I(signal_light_c), .O(signal_light));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[14:26])
    OB expansion3_pad (.I(expansion3_c_11), .O(expansion3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    OB expansion2_pad (.I(expansion2_c_10), .O(expansion2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    OB expansion1_pad (.I(expansion1_c_9), .O(expansion1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[14:24])
    OB Stepper_A_En_pad (.I(Stepper_A_En_c), .O(Stepper_A_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    LUT4 Select_4283_i2_2_lut_3_lut_4_lut (.A(n32261), .B(n32168), .C(read_value_adj_1055[3]), 
         .D(rw), .Z(n2_adj_925)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4283_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4284_i2_2_lut_3_lut_4_lut (.A(n32261), .B(n32168), .C(read_value_adj_1055[2]), 
         .D(rw), .Z(n2_adj_929)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4284_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4280_i2_2_lut_3_lut_4_lut (.A(n32261), .B(n32168), .C(read_value_adj_1055[6]), 
         .D(rw), .Z(n2_adj_919)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4280_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    OB Stepper_A_M2_pad (.I(Stepper_A_M2_c_2), .O(Stepper_A_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    OB Stepper_A_M1_pad (.I(Stepper_A_M1_c_1), .O(Stepper_A_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    LUT4 i1_2_lut_rep_338_3_lut_4_lut (.A(n32233), .B(n32251), .C(rw), 
         .D(prev_select_adj_634), .Z(n32159)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_338_3_lut_4_lut.init = 16'h0004;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(n32233), .B(n32251), .C(n34065), 
         .D(prev_select_adj_634), .Z(n2769)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i23207_4_lut_rep_501 (.A(reset_count[14]), .B(n205), .C(n29544), 
         .D(n29953), .Z(n34067)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23207_4_lut_rep_501.init = 16'h575f;
    LUT4 i15_2_lut_rep_343_3_lut_4_lut (.A(register_addr[4]), .B(n32234), 
         .C(n34064), .D(select[3]), .Z(n32164)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam i15_2_lut_rep_343_3_lut_4_lut.init = 16'h2000;
    LUT4 i114_2_lut_3_lut_4_lut (.A(register_addr[4]), .B(n32234), .C(prev_select_adj_881), 
         .D(select[3]), .Z(n178)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam i114_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 Select_4297_i9_2_lut_3_lut_4_lut (.A(register_addr[4]), .B(n32234), 
         .C(read_size_adj_1101[0]), .D(select[3]), .Z(n9_adj_923)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4297_i9_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i15_2_lut_rep_340_3_lut_4_lut (.A(register_addr[4]), .B(n32234), 
         .C(rw), .D(select[3]), .Z(n32161)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam i15_2_lut_rep_340_3_lut_4_lut.init = 16'hd000;
    LUT4 i114_2_lut_3_lut_4_lut_adj_482 (.A(register_addr[4]), .B(n32234), 
         .C(prev_select_adj_844), .D(select[3]), .Z(n14271)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam i114_2_lut_3_lut_4_lut_adj_482.init = 16'h0d00;
    LUT4 i23207_4_lut_rep_499 (.A(reset_count[14]), .B(n205), .C(n29544), 
         .D(n29953), .Z(n34065)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23207_4_lut_rep_499.init = 16'h575f;
    LUT4 i23207_4_lut_rep_504 (.A(reset_count[14]), .B(n205), .C(n29544), 
         .D(n29953), .Z(n34070)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23207_4_lut_rep_504.init = 16'h575f;
    LUT4 i23207_4_lut_rep_505 (.A(reset_count[14]), .B(n205), .C(n29544), 
         .D(n29953), .Z(n34071)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23207_4_lut_rep_505.init = 16'h575f;
    LUT4 Select_4266_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[12]), 
         .D(rw), .Z(n2_adj_569)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4266_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4278_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[8]), 
         .D(n34064), .Z(n2_adj_845)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4278_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4275_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[9]), 
         .D(rw), .Z(n2_adj_635)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4275_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4272_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[10]), 
         .D(rw), .Z(n2_adj_809)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4272_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4269_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[11]), 
         .D(rw), .Z(n2_adj_584)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4269_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_adj_483 (.A(n32252), .B(n32251), .C(n34065), 
         .D(prev_select_adj_722), .Z(n13476)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut_adj_483.init = 16'h0008;
    LUT4 i1_2_lut_rep_344_3_lut_4_lut (.A(n32252), .B(n32251), .C(rw), 
         .D(prev_select_adj_722), .Z(n32165)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_344_3_lut_4_lut.init = 16'h0008;
    LUT4 Select_4279_i3_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[7]), 
         .D(n34064), .Z(n3)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4279_i3_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4280_i3_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[6]), 
         .D(rw), .Z(n3_adj_900)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4280_i3_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i30_2_lut_rep_469 (.A(uart_rx_c), .B(prev_uart_rx), .Z(n32290)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(475[7:30])
    defparam i30_2_lut_rep_469.init = 16'h2222;
    LUT4 Select_4281_i3_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[5]), 
         .D(rw), .Z(n3_adj_906)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4281_i3_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2737_2_lut_3_lut (.A(uart_rx_c), .B(prev_uart_rx), .C(n7787), 
         .Z(n14355)) /* synthesis lut_function=(!(A (B (C))+!A (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(475[7:30])
    defparam i2737_2_lut_3_lut.init = 16'h2f2f;
    LUT4 i15832_2_lut_3_lut (.A(uart_rx_c), .B(prev_uart_rx), .C(n658[0]), 
         .Z(n99_adj_1349[0])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(475[7:30])
    defparam i15832_2_lut_3_lut.init = 16'hd0d0;
    LUT4 Select_4282_i3_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[4]), 
         .D(rw), .Z(n3_adj_882)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4282_i3_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4283_i3_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[3]), 
         .D(rw), .Z(n3_adj_924)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4283_i3_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4284_i3_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[2]), 
         .D(rw), .Z(n3_adj_928)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4284_i3_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4285_i3_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[1]), 
         .D(rw), .Z(n3_adj_931)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4285_i3_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1P3AX reset_count_2657_2658__i1 (.D(n66_adj_1469[0]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658__i1.GSR = "ENABLED";
    LUT4 Select_4263_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[13]), 
         .D(rw), .Z(n2_adj_724)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4263_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i23166_2_lut (.A(n30566), .B(n34065), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23166_2_lut.init = 16'heeee;
    LUT4 Select_4286_i3_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[0]), 
         .D(rw), .Z(n3_adj_926)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4286_i3_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4209_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[31]), 
         .D(rw), .Z(n2_adj_598)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4209_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4212_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[30]), 
         .D(rw), .Z(n2_adj_579)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4212_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4215_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[29]), 
         .D(rw), .Z(n2_adj_904)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4215_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i23164_4_lut (.A(reset_count[0]), .B(n142), .C(n10), .D(n29544), 
         .Z(n30566)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i23164_4_lut.init = 16'h0001;
    LUT4 Select_4218_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[28]), 
         .D(rw), .Z(n2_adj_725)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4218_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4221_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[27]), 
         .D(rw), .Z(n2_adj_903)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4221_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4224_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[26]), 
         .D(rw), .Z(n2_adj_597)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4224_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i4_4_lut (.A(reset_count[5]), .B(reset_count[1]), .C(reset_count[2]), 
         .D(reset_count[3]), .Z(n10)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(458[13:24])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 Select_4227_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[25]), 
         .D(rw), .Z(n2_adj_681)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4227_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4230_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[24]), 
         .D(rw), .Z(n2_adj_637)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4230_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4233_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[23]), 
         .D(rw), .Z(n2_adj_583)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4233_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4236_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[22]), 
         .D(rw), .Z(n2_adj_808)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4236_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4239_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[21]), 
         .D(rw), .Z(n2)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4239_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut (.A(reset_count[7]), .B(reset_count[8]), .Z(n142)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(458[13:24])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 Select_4242_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[20]), 
         .D(rw), .Z(n2_adj_677)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4242_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4245_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[19]), 
         .D(rw), .Z(n2_adj_933)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4245_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4248_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[18]), 
         .D(rw), .Z(n2_adj_806)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4248_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4251_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[17]), 
         .D(rw), .Z(n2_adj_580)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4251_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4254_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[16]), 
         .D(rw), .Z(n2_adj_586)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4254_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4257_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[15]), 
         .D(rw), .Z(n2_adj_901)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4257_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_4260_i2_2_lut_3_lut_4_lut (.A(n32252), .B(n32251), .C(read_value_adj_1017[14]), 
         .D(rw), .Z(n2_adj_897)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_4260_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_3_lut (.A(reset_count[12]), .B(reset_count[11]), .C(reset_count[13]), 
         .Z(n29544)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(458[13:24])
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i23207_4_lut_rep_395 (.A(reset_count[14]), .B(n205), .C(n29544), 
         .D(n29953), .Z(n32216)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23207_4_lut_rep_395.init = 16'h575f;
    LUT4 i1_2_lut_4_lut (.A(count_adj_1267[4]), .B(count_adj_1267[3]), .C(n32257), 
         .D(n29947), .Z(n29948)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfe00;
    LUT4 i23207_4_lut_rep_500 (.A(reset_count[14]), .B(n205), .C(n29544), 
         .D(n29953), .Z(n34066)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23207_4_lut_rep_500.init = 16'h575f;
    LUT4 i23207_4_lut_rep_502 (.A(reset_count[14]), .B(n205), .C(n29544), 
         .D(n29953), .Z(n34068)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23207_4_lut_rep_502.init = 16'h575f;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32172), .B(n32306), .C(register_addr[0]), 
         .D(n34065), .Z(n11961)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[17:42])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf040;
    LUT4 i23215_4_lut (.A(n32294), .B(n32296), .C(n28329), .D(n28144), 
         .Z(n30617)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;
    defparam i23215_4_lut.init = 16'h5455;
    LUT4 i2_3_lut_rep_481 (.A(count_adj_1267[2]), .B(count_adj_1267[3]), 
         .C(count_adj_1267[1]), .Z(n32302)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_rep_481.init = 16'h8080;
    LUT4 i1_2_lut_rep_424_4_lut (.A(count_adj_1267[2]), .B(count_adj_1267[3]), 
         .C(count_adj_1267[1]), .D(count_adj_1267[0]), .Z(n32245)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_424_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_484 (.A(n32172), .B(n32306), .C(register_addr[0]), 
         .D(n34065), .Z(n13598)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C)+!B (C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[17:42])
    defparam i1_2_lut_3_lut_4_lut_adj_484.init = 16'h0f04;
    LUT4 i1_2_lut_rep_485 (.A(select[5]), .B(prev_select_adj_893), .Z(n32306)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[17:42])
    defparam i1_2_lut_rep_485.init = 16'h2222;
    LUT4 i1_2_lut_rep_341_2_lut_3_lut (.A(select[5]), .B(prev_select_adj_893), 
         .C(n34065), .Z(n32162)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[17:42])
    defparam i1_2_lut_rep_341_2_lut_3_lut.init = 16'h0202;
    LUT4 n44_bdd_4_lut (.A(n44_adj_575), .B(n30320), .C(count_adj_1215[9]), 
         .D(n30308), .Z(n32125)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n44_bdd_4_lut.init = 16'h00ca;
    OB Stepper_A_M0_pad (.I(Stepper_A_M0_c_0), .O(Stepper_A_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:29])
    LUT4 i1_4_lut (.A(n34065), .B(state_adj_1287[2]), .C(state_adj_1287[3]), 
         .D(n29883), .Z(n29194)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[17:42])
    defparam i1_4_lut.init = 16'h1410;
    LUT4 i1_2_lut_adj_485 (.A(state_adj_1287[1]), .B(state_adj_1287[0]), 
         .Z(n29883)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[17:42])
    defparam i1_2_lut_adj_485.init = 16'h8888;
    LUT4 i2_4_lut (.A(n29953), .B(n28017), .C(reset_count[11]), .D(reset_count[8]), 
         .Z(n29954)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'ha080;
    LUT4 i2_3_lut_adj_486 (.A(reset_count[6]), .B(reset_count[5]), .C(reset_count[7]), 
         .Z(n28017)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(458[13:24])
    defparam i2_3_lut_adj_486.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_487 (.A(count_adj_1267[0]), .B(n32302), 
         .C(n32258), .D(n32256), .Z(n30001)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_487.init = 16'h8000;
    LUT4 i1_2_lut_adj_488 (.A(reset_count[10]), .B(reset_count[9]), .Z(n29953)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_488.init = 16'h8888;
    LUT4 i3_4_lut_4_lut (.A(n34065), .B(n32282), .C(n32315), .D(n29920), 
         .Z(n13118)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i3_4_lut_4_lut.init = 16'h0100;
    LUT4 i15812_2_lut_2_lut (.A(n34065), .B(databus[7]), .Z(n281[15])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i15812_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_rep_368_3_lut_4_lut (.A(select[4]), .B(n32315), .C(prev_select_adj_722), 
         .D(n32252), .Z(n32189)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_rep_368_3_lut_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_rep_382_3_lut_4_lut (.A(select[4]), .B(n32315), .C(n32279), 
         .D(n32282), .Z(n32203)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_rep_382_3_lut_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_rep_394_3_lut_4_lut (.A(register_addr[5]), .B(n32316), 
         .C(n32315), .D(select[4]), .Z(n32215)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_rep_394_3_lut_4_lut.init = 16'h0200;
    LUT4 i2_3_lut_rep_336_4_lut (.A(select[3]), .B(n32205), .C(n32235), 
         .D(prev_select_adj_881), .Z(n32157)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam i2_3_lut_rep_336_4_lut.init = 16'h0080;
    LUT4 Select_4285_i10_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1100[1]), 
         .D(n34064), .Z(n10_adj_930)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4285_i10_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i23219_4_lut (.A(n32264), .B(n5_adj_912), .C(n28330), .D(n28132), 
         .Z(n30621)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i23219_4_lut.init = 16'h3233;
    LUT4 i23145_4_lut (.A(n30546), .B(n17), .C(n15), .D(n16), .Z(n28407)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i23145_4_lut.init = 16'h8000;
    LUT4 i23144_4_lut (.A(n29), .B(n42), .C(n38), .D(n30_adj_899), .Z(n30546)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i23144_4_lut.init = 16'h0001;
    LUT4 n44_bdd_4_lut_adj_489 (.A(n44_adj_726), .B(n30324), .C(count_adj_1228[9]), 
         .D(n30302), .Z(n32127)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n44_bdd_4_lut_adj_489.init = 16'h00ca;
    LUT4 i7_4_lut (.A(timeout_count[16]), .B(timeout_count[25]), .C(timeout_count[15]), 
         .D(timeout_count[24]), .Z(n17)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i15080_2_lut_2_lut (.A(n34065), .B(n8447), .Z(n107)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i15080_2_lut_2_lut.init = 16'h4444;
    FD1P3IX timeout_count__i31 (.D(n658[31]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i31.GSR = "ENABLED";
    LUT4 i5_2_lut (.A(timeout_count[8]), .B(timeout_count[20]), .Z(n15)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5_2_lut.init = 16'h8888;
    LUT4 i15256_2_lut_2_lut (.A(n34065), .B(databus[2]), .Z(n580_adj_1036[2])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i15256_2_lut_2_lut.init = 16'h4444;
    LUT4 i15395_2_lut_2_lut (.A(n34065), .B(databus[4]), .Z(n580_adj_998[4])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i15395_2_lut_2_lut.init = 16'h4444;
    LUT4 i6_4_lut (.A(timeout_count[17]), .B(timeout_count[9]), .C(timeout_count[23]), 
         .D(timeout_count[10]), .Z(n16)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_331_3_lut_4_lut (.A(select[4]), .B(n32199), .C(prev_select_adj_773), 
         .D(n32261), .Z(n32152)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_rep_331_3_lut_4_lut.init = 16'h0200;
    LUT4 i7_2_lut (.A(timeout_count[5]), .B(timeout_count[18]), .Z(n29)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 Select_4269_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[11]), 
         .D(rw), .Z(n8_adj_683)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4269_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4266_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[12]), 
         .D(rw), .Z(n8_adj_570)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4266_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_3_lut_rep_339_4_lut (.A(select[3]), .B(n32205), .C(n32204), 
         .D(prev_select_adj_844), .Z(n32160)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam i2_3_lut_rep_339_4_lut.init = 16'h0020;
    FD1P3IX timeout_count__i30 (.D(n658[30]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i30.GSR = "ENABLED";
    FD1P3IX timeout_count__i29 (.D(n658[29]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i29.GSR = "ENABLED";
    FD1P3IX timeout_count__i28 (.D(n658[28]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i28.GSR = "ENABLED";
    FD1P3IX timeout_count__i27 (.D(n658[27]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i27.GSR = "ENABLED";
    FD1P3IX timeout_count__i26 (.D(n658[26]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i26.GSR = "ENABLED";
    FD1P3IX timeout_count__i25 (.D(n658[25]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i25.GSR = "ENABLED";
    FD1P3IX timeout_count__i24 (.D(n658[24]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i24.GSR = "ENABLED";
    FD1P3IX timeout_count__i23 (.D(n658[23]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i23.GSR = "ENABLED";
    FD1P3IX timeout_count__i22 (.D(n658[22]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i22.GSR = "ENABLED";
    FD1P3IX timeout_count__i21 (.D(n658[21]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i21.GSR = "ENABLED";
    LUT4 i20_4_lut (.A(timeout_count[12]), .B(n40), .C(n34_adj_898), .D(timeout_count[19]), 
         .Z(n42)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i23213_4_lut (.A(n32317), .B(n32283), .C(n28331), .D(n28133), 
         .Z(n30615)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i23213_4_lut.init = 16'h3233;
    FD1P3IX timeout_count__i20 (.D(n658[20]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i20.GSR = "ENABLED";
    FD1P3IX timeout_count__i19 (.D(n658[19]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i19.GSR = "ENABLED";
    FD1P3IX timeout_count__i18 (.D(n658[18]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i18.GSR = "ENABLED";
    FD1P3IX timeout_count__i17 (.D(n658[17]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i17.GSR = "ENABLED";
    FD1P3IX timeout_count__i16 (.D(n658[16]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i16.GSR = "ENABLED";
    FD1P3IX timeout_count__i15 (.D(n658[15]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i15.GSR = "ENABLED";
    FD1P3IX timeout_count__i14 (.D(n658[14]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i14.GSR = "ENABLED";
    FD1P3IX timeout_count__i13 (.D(n658[13]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i13.GSR = "ENABLED";
    FD1P3IX timeout_count__i12 (.D(n658[12]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i12.GSR = "ENABLED";
    FD1P3IX timeout_count__i11 (.D(n658[11]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i11.GSR = "ENABLED";
    FD1P3IX timeout_count__i10 (.D(n658[10]), .SP(n9309), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i10.GSR = "ENABLED";
    FD1P3IX timeout_count__i9 (.D(n658[9]), .SP(n14355), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i9.GSR = "ENABLED";
    FD1P3IX timeout_count__i8 (.D(n658[8]), .SP(n14355), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i8.GSR = "ENABLED";
    FD1P3IX timeout_count__i7 (.D(n658[7]), .SP(n14355), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i7.GSR = "ENABLED";
    FD1P3IX timeout_count__i6 (.D(n658[6]), .SP(n14355), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i6.GSR = "ENABLED";
    FD1P3IX timeout_count__i5 (.D(n658[5]), .SP(n14355), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i5.GSR = "ENABLED";
    FD1P3IX timeout_count__i4 (.D(n658[4]), .SP(n14355), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i4.GSR = "ENABLED";
    FD1P3IX timeout_count__i3 (.D(n658[3]), .SP(n14355), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i3.GSR = "ENABLED";
    FD1P3IX timeout_count__i2 (.D(n658[2]), .SP(n14355), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i2.GSR = "ENABLED";
    FD1P3IX timeout_count__i1 (.D(n658[1]), .SP(n14355), .CD(n32290), 
            .CK(debug_c_c), .Q(timeout_count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(472[9] 490[6])
    defparam timeout_count__i1.GSR = "ENABLED";
    LUT4 i16_4_lut (.A(timeout_count[31]), .B(timeout_count[22]), .C(timeout_count[21]), 
         .D(timeout_count[28]), .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_4_lut (.A(n34065), .B(n32261), .C(n32199), .D(n32152), 
         .Z(n9496)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (D)))) */ ;
    defparam i2_4_lut_4_lut.init = 16'h5100;
    LUT4 Select_4272_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[10]), 
         .D(n34064), .Z(n8_adj_846)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4272_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4275_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[9]), 
         .D(rw), .Z(n8_adj_727)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4275_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    OB Stepper_A_Dir_pad (.I(Stepper_A_Dir_c), .O(Stepper_A_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:30])
    OB Stepper_A_Step_pad (.I(Stepper_A_Step_c), .O(Stepper_A_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(392[17:31])
    OB Stepper_Z_En_pad (.I(Stepper_Z_En_c), .O(Stepper_Z_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    OB Stepper_Z_M2_pad (.I(Stepper_Z_M2_c_2), .O(Stepper_Z_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    OB Stepper_Z_M1_pad (.I(Stepper_Z_M1_c_1), .O(Stepper_Z_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    OB Stepper_Z_M0_pad (.I(Stepper_Z_M0_c_0), .O(Stepper_Z_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:29])
    OB Stepper_Z_Dir_pad (.I(Stepper_Z_Dir_c), .O(Stepper_Z_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:30])
    OB Stepper_Z_Step_pad (.I(Stepper_Z_Step_c), .O(Stepper_Z_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(384[17:31])
    OB Stepper_Y_En_pad (.I(Stepper_Y_En_c), .O(Stepper_Y_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    OB Stepper_Y_M2_pad (.I(Stepper_Y_M2_c_2), .O(Stepper_Y_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    OB Stepper_Y_M1_pad (.I(Stepper_Y_M1_c_1), .O(Stepper_Y_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    OB Stepper_Y_M0_pad (.I(Stepper_Y_M0_c_0), .O(Stepper_Y_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:29])
    OB Stepper_Y_Dir_pad (.I(Stepper_Y_Dir_c), .O(Stepper_Y_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:30])
    OB Stepper_Y_Step_pad (.I(Stepper_Y_Step_c), .O(Stepper_Y_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(376[17:31])
    OB Stepper_X_En_pad (.I(Stepper_X_En_c), .O(Stepper_X_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    OB Stepper_X_M2_pad (.I(Stepper_X_M2_c_2), .O(Stepper_X_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    OB Stepper_X_M1_pad (.I(Stepper_X_M1_c_1), .O(Stepper_X_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    OB Stepper_X_M0_pad (.I(Stepper_X_M0_c_0), .O(Stepper_X_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:29])
    OB Stepper_X_Dir_pad (.I(Stepper_X_Dir_c), .O(Stepper_X_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:30])
    OB Stepper_X_Step_pad (.I(Stepper_X_Step_c), .O(Stepper_X_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(368[17:31])
    OB status_led_pad_0 (.I(VCC_net), .O(status_led[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    OB status_led_pad_1 (.I(VCC_net), .O(status_led[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    OB status_led_pad_2 (.I(VCC_net), .O(status_led[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[20:30])
    OB uart_tx_pad (.I(uart_tx_c), .O(uart_tx));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[14:21])
    BB expansion4_pad (.I(n10948), .T(n10947), .B(expansion4), .O(expansion4_out));
    LUT4 i1_2_lut_rep_333_3_lut_4_lut (.A(select[4]), .B(n32199), .C(prev_select_adj_675), 
         .D(n32305), .Z(n32154)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_rep_333_3_lut_4_lut.init = 16'h0200;
    LUT4 Select_4278_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[8]), 
         .D(rw), .Z(n8_adj_680)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4278_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i20_2_lut_3_lut_4_lut (.A(select[4]), .B(n32199), .C(rw), .D(n32305), 
         .Z(n52_adj_676)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i20_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4263_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[13]), 
         .D(n34064), .Z(n8_adj_573)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4263_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4209_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[31]), 
         .D(rw), .Z(n8_adj_918)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4209_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4212_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[30]), 
         .D(n34064), .Z(n8_adj_568)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4212_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4215_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[29]), 
         .D(rw), .Z(n8_adj_922)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4215_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    CCU2D add_20289_24 (.A0(timeout_count[31]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(battery_voltage[15]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27737), .S1(n7787));
    defparam add_20289_24.INIT0 = 16'h5555;
    defparam add_20289_24.INIT1 = 16'h0000;
    defparam add_20289_24.INJECT1_0 = "NO";
    defparam add_20289_24.INJECT1_1 = "NO";
    CCU2D add_20289_22 (.A0(timeout_count[29]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[30]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27736), .COUT(n27737));
    defparam add_20289_22.INIT0 = 16'h5555;
    defparam add_20289_22.INIT1 = 16'h5555;
    defparam add_20289_22.INJECT1_0 = "NO";
    defparam add_20289_22.INJECT1_1 = "NO";
    CCU2D add_20289_20 (.A0(timeout_count[27]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[28]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27735), .COUT(n27736));
    defparam add_20289_20.INIT0 = 16'h5555;
    defparam add_20289_20.INIT1 = 16'h5555;
    defparam add_20289_20.INJECT1_0 = "NO";
    defparam add_20289_20.INJECT1_1 = "NO";
    CCU2D add_20289_18 (.A0(timeout_count[25]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[26]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27734), .COUT(n27735));
    defparam add_20289_18.INIT0 = 16'h5aaa;
    defparam add_20289_18.INIT1 = 16'h5555;
    defparam add_20289_18.INJECT1_0 = "NO";
    defparam add_20289_18.INJECT1_1 = "NO";
    CCU2D add_20289_16 (.A0(timeout_count[23]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[24]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27733), .COUT(n27734));
    defparam add_20289_16.INIT0 = 16'h5aaa;
    defparam add_20289_16.INIT1 = 16'h5aaa;
    defparam add_20289_16.INJECT1_0 = "NO";
    defparam add_20289_16.INJECT1_1 = "NO";
    CCU2D add_31_33 (.A0(timeout_count[31]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(battery_voltage[15]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27046), 
          .S0(n658[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_33.INIT0 = 16'h5aaa;
    defparam add_31_33.INIT1 = 16'h0000;
    defparam add_31_33.INJECT1_0 = "NO";
    defparam add_31_33.INJECT1_1 = "NO";
    CCU2D add_31_31 (.A0(timeout_count[29]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[30]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27045), 
          .COUT(n27046), .S0(n658[29]), .S1(n658[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_31.INIT0 = 16'h5aaa;
    defparam add_31_31.INIT1 = 16'h5aaa;
    defparam add_31_31.INJECT1_0 = "NO";
    defparam add_31_31.INJECT1_1 = "NO";
    CCU2D add_20289_14 (.A0(timeout_count[21]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[22]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27732), .COUT(n27733));
    defparam add_20289_14.INIT0 = 16'h5555;
    defparam add_20289_14.INIT1 = 16'h5555;
    defparam add_20289_14.INJECT1_0 = "NO";
    defparam add_20289_14.INJECT1_1 = "NO";
    CCU2D add_31_13 (.A0(timeout_count[11]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[12]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27036), 
          .COUT(n27037), .S0(n658[11]), .S1(n658[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_13.INIT0 = 16'h5aaa;
    defparam add_31_13.INIT1 = 16'h5aaa;
    defparam add_31_13.INJECT1_0 = "NO";
    defparam add_31_13.INJECT1_1 = "NO";
    CCU2D add_31_11 (.A0(timeout_count[9]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[10]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27035), 
          .COUT(n27036), .S0(n658[9]), .S1(n658[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_11.INIT0 = 16'h5aaa;
    defparam add_31_11.INIT1 = 16'h5aaa;
    defparam add_31_11.INJECT1_0 = "NO";
    defparam add_31_11.INJECT1_1 = "NO";
    CCU2D add_20289_12 (.A0(timeout_count[19]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[20]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27731), .COUT(n27732));
    defparam add_20289_12.INIT0 = 16'h5555;
    defparam add_20289_12.INIT1 = 16'h5aaa;
    defparam add_20289_12.INJECT1_0 = "NO";
    defparam add_20289_12.INJECT1_1 = "NO";
    CCU2D add_20289_10 (.A0(timeout_count[17]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[18]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27730), .COUT(n27731));
    defparam add_20289_10.INIT0 = 16'h5aaa;
    defparam add_20289_10.INIT1 = 16'h5555;
    defparam add_20289_10.INJECT1_0 = "NO";
    defparam add_20289_10.INJECT1_1 = "NO";
    CCU2D add_20289_8 (.A0(timeout_count[15]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[16]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27729), .COUT(n27730));
    defparam add_20289_8.INIT0 = 16'h5aaa;
    defparam add_20289_8.INIT1 = 16'h5aaa;
    defparam add_20289_8.INJECT1_0 = "NO";
    defparam add_20289_8.INJECT1_1 = "NO";
    CCU2D add_20289_6 (.A0(timeout_count[13]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[14]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27728), .COUT(n27729));
    defparam add_20289_6.INIT0 = 16'h5555;
    defparam add_20289_6.INIT1 = 16'h5555;
    defparam add_20289_6.INJECT1_0 = "NO";
    defparam add_20289_6.INJECT1_1 = "NO";
    LUT4 Select_4218_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[28]), 
         .D(rw), .Z(n8_adj_907)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4218_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4221_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[27]), 
         .D(rw), .Z(n8_adj_585)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4221_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4224_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[26]), 
         .D(rw), .Z(n8_adj_921)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4224_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4227_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[25]), 
         .D(rw), .Z(n8_adj_679)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4227_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4297_i5_2_lut_3_lut_4_lut (.A(select[4]), .B(n32199), .C(read_size_adj_980[0]), 
         .D(n32305), .Z(n5)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam Select_4297_i5_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4230_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[24]), 
         .D(n34064), .Z(n8_adj_684)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4230_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4233_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[23]), 
         .D(rw), .Z(n8_adj_678)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4233_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    FD1P3AX reset_count_2657_2658__i2 (.D(n66_adj_1469[1]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658__i2.GSR = "ENABLED";
    LUT4 Select_4236_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[22]), 
         .D(rw), .Z(n8)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4236_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    CCU2D add_20289_4 (.A0(timeout_count[11]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(timeout_count[12]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27727), .COUT(n27728));
    defparam add_20289_4.INIT0 = 16'h5555;
    defparam add_20289_4.INIT1 = 16'h5555;
    defparam add_20289_4.INJECT1_0 = "NO";
    defparam add_20289_4.INJECT1_1 = "NO";
    CCU2D add_20289_2 (.A0(timeout_count[9]), .B0(timeout_count[8]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[10]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .COUT(n27727));
    defparam add_20289_2.INIT0 = 16'h7000;
    defparam add_20289_2.INIT1 = 16'h5aaa;
    defparam add_20289_2.INJECT1_0 = "NO";
    defparam add_20289_2.INJECT1_1 = "NO";
    LUT4 Select_4239_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[21]), 
         .D(n34064), .Z(n8_adj_682)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4239_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4242_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[20]), 
         .D(n34064), .Z(n8_adj_934)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4242_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4245_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[19]), 
         .D(n34064), .Z(n8_adj_932)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4245_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4248_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[18]), 
         .D(n34064), .Z(n8_adj_636)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4248_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4251_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[17]), 
         .D(n34064), .Z(n8_adj_902)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4251_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    CCU2D add_31_29 (.A0(timeout_count[27]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[28]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27044), 
          .COUT(n27045), .S0(n658[27]), .S1(n658[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_29.INIT0 = 16'h5aaa;
    defparam add_31_29.INIT1 = 16'h5aaa;
    defparam add_31_29.INJECT1_0 = "NO";
    defparam add_31_29.INJECT1_1 = "NO";
    CCU2D add_31_27 (.A0(timeout_count[25]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[26]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27043), 
          .COUT(n27044), .S0(n658[25]), .S1(n658[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_27.INIT0 = 16'h5aaa;
    defparam add_31_27.INIT1 = 16'h5aaa;
    defparam add_31_27.INJECT1_0 = "NO";
    defparam add_31_27.INJECT1_1 = "NO";
    LUT4 Select_4254_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[16]), 
         .D(n34064), .Z(n8_adj_582)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4254_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4257_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[15]), 
         .D(n34064), .Z(n8_adj_578)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4257_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_4260_i8_2_lut_3_lut_4_lut (.A(select[3]), .B(n32205), .C(read_value_adj_1092[14]), 
         .D(n34064), .Z(n8_adj_896)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(653[4] 669[11])
    defparam Select_4260_i8_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i23207_4_lut_rep_503 (.A(reset_count[14]), .B(n205), .C(n29544), 
         .D(n29953), .Z(n34069)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i23207_4_lut_rep_503.init = 16'h575f;
    FD1P3AX reset_count_2657_2658__i3 (.D(n66_adj_1469[2]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658__i3.GSR = "ENABLED";
    FD1P3AX reset_count_2657_2658__i4 (.D(n66_adj_1469[3]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658__i4.GSR = "ENABLED";
    FD1P3AX reset_count_2657_2658__i5 (.D(n66_adj_1469[4]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658__i5.GSR = "ENABLED";
    FD1P3AX reset_count_2657_2658__i6 (.D(n66_adj_1469[5]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658__i6.GSR = "ENABLED";
    FD1P3AX reset_count_2657_2658__i7 (.D(n66_adj_1469[6]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658__i7.GSR = "ENABLED";
    FD1P3AX reset_count_2657_2658__i8 (.D(n66_adj_1469[7]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658__i8.GSR = "ENABLED";
    FD1P3AX reset_count_2657_2658__i9 (.D(n66_adj_1469[8]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658__i9.GSR = "ENABLED";
    FD1P3AX reset_count_2657_2658__i10 (.D(n66_adj_1469[9]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658__i10.GSR = "ENABLED";
    FD1P3AX reset_count_2657_2658__i11 (.D(n66_adj_1469[10]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658__i11.GSR = "ENABLED";
    FD1P3AX reset_count_2657_2658__i12 (.D(n66_adj_1469[11]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658__i12.GSR = "ENABLED";
    FD1P3AX reset_count_2657_2658__i13 (.D(n66_adj_1469[12]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658__i13.GSR = "ENABLED";
    FD1P3AX reset_count_2657_2658__i14 (.D(n66_adj_1469[13]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658__i14.GSR = "ENABLED";
    FD1P3AX reset_count_2657_2658__i15 (.D(n66_adj_1469[14]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658__i15.GSR = "ENABLED";
    GSR GSR_INST (.GSR(VCC_net));
    LUT4 n44_bdd_4_lut_adj_490 (.A(n44), .B(n30330), .C(count_adj_1267[9]), 
         .D(n30304), .Z(n32129)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n44_bdd_4_lut_adj_490.init = 16'h00ca;
    CCU2D add_31_25 (.A0(timeout_count[23]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[24]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27042), 
          .COUT(n27043), .S0(n658[23]), .S1(n658[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_25.INIT0 = 16'h5aaa;
    defparam add_31_25.INIT1 = 16'h5aaa;
    defparam add_31_25.INJECT1_0 = "NO";
    defparam add_31_25.INJECT1_1 = "NO";
    LUT4 i9997_3_lut_4_lut_4_lut (.A(n34065), .B(n32204), .C(n32187), 
         .D(n32306), .Z(n16718)) /* synthesis lut_function=(!(A+!(B (D)+!B !(C+!(D))))) */ ;
    defparam i9997_3_lut_4_lut_4_lut.init = 16'h4500;
    LUT4 i2_3_lut_4_lut_4_lut (.A(n34065), .B(n32200), .C(prev_select_adj_634), 
         .D(n32203), .Z(n9485)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_4_lut_4_lut.init = 16'h0400;
    CCU2D add_31_23 (.A0(timeout_count[21]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[22]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27041), 
          .COUT(n27042), .S0(n658[21]), .S1(n658[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_23.INIT0 = 16'h5aaa;
    defparam add_31_23.INIT1 = 16'h5aaa;
    defparam add_31_23.INJECT1_0 = "NO";
    defparam add_31_23.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_491 (.A(div_factor_reg_adj_1015[9]), .B(register_addr[1]), 
         .C(steps_reg_adj_1016[9]), .D(register_addr[0]), .Z(n29860)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_4_lut_adj_491.init = 16'hc088;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n34065), .B(prev_select_adj_773), 
         .C(n32168), .D(n32261), .Z(n14114)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h1000;
    LUT4 i1_4_lut_adj_492 (.A(count_adj_1215[8]), .B(n32293), .C(count_adj_1215[5]), 
         .D(n41), .Z(n44_adj_575)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_adj_492.init = 16'heaaa;
    LUT4 i23154_3_lut (.A(count_adj_1215[8]), .B(count_adj_1215[6]), .C(n5_adj_920), 
         .Z(n30320)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i23154_3_lut.init = 16'h0101;
    LUT4 i14764_3_lut (.A(Stepper_A_Dir_c), .B(div_factor_reg_adj_1053[5]), 
         .C(register_addr[1]), .Z(n21453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i14764_3_lut.init = 16'hcaca;
    \ArmPeripheral(axis_haddr=8'b0100000)  arm_z (.limit_c_2(limit_c_2), .Stepper_Z_M0_c_0(Stepper_Z_M0_c_0), 
            .register_addr({register_addr}), .debug_c_c(debug_c_c), .VCC_net(VCC_net), 
            .GND_net(battery_voltage[15]), .Stepper_Z_nFault_c(Stepper_Z_nFault_c), 
            .n34066(n34066), .n3948({n3948}), .\read_size[0] (read_size_adj_1018[0]), 
            .n13476(n13476), .n28302(n28302), .n579(n571[0]), .prev_step_clk(prev_step_clk_adj_687), 
            .step_clk(step_clk_adj_686), .n13769(n13769), .prev_select(prev_select_adj_722), 
            .n32215(n32215), .n34067(n34067), .\databus[31] (databus[31]), 
            .\databus[30] (databus[30]), .\databus[29] (databus[29]), .\databus[28] (databus[28]), 
            .\databus[27] (databus[27]), .\databus[26] (databus[26]), .\databus[25] (databus[25]), 
            .\databus[24] (databus[24]), .\databus[23] (databus[23]), .\databus[22] (databus[22]), 
            .\databus[21] (databus[21]), .\databus[20] (databus[20]), .\databus[19] (databus[19]), 
            .\databus[18] (databus[18]), .\databus[17] (databus[17]), .\databus[16] (databus[16]), 
            .\databus[15] (databus[15]), .n34068(n34068), .\databus[13] (databus[13]), 
            .\databus[11] (databus[11]), .\databus[10] (databus[10]), .\div_factor_reg[9] (div_factor_reg_adj_1015[9]), 
            .\databus[9] (databus[9]), .\databus[7] (databus[7]), .\div_factor_reg[6] (div_factor_reg_adj_1015[6]), 
            .\databus[6] (databus[6]), .\div_factor_reg[5] (div_factor_reg_adj_1015[5]), 
            .\databus[5] (databus[5]), .n608(n580_adj_998[4]), .n610(n580_adj_1036[2]), 
            .\control_reg[7] (control_reg_adj_1014[7]), .Stepper_Z_En_c(Stepper_Z_En_c), 
            .Stepper_Z_Dir_c(Stepper_Z_Dir_c), .\control_reg[3] (control_reg_adj_1014[3]), 
            .\databus[3] (databus[3]), .Stepper_Z_M2_c_2(Stepper_Z_M2_c_2), 
            .Stepper_Z_M1_c_1(Stepper_Z_M1_c_1), .\databus[1] (databus[1]), 
            .\read_size[2] (read_size_adj_1018[2]), .n30020(n30020), .n34070(n34070), 
            .\steps_reg[9] (steps_reg_adj_1016[9]), .\steps_reg[6] (steps_reg_adj_1016[6]), 
            .n34071(n34071), .\steps_reg[5] (steps_reg_adj_1016[5]), .\steps_reg[3] (steps_reg_adj_1016[3]), 
            .n32315(n32315), .n29750(n29750), .n32232(n32232), .n32234(n32234), 
            .n32316(n32316), .n32200(n32200), .n32205(n32205), .\select[4] (select[4]), 
            .n32251(n32251), .n32253(n32253), .rw(rw), .n32189(n32189), 
            .n32252(n32252), .n32199(n32199), .n32166(n32166), .n32314(n32314), 
            .n9(n9), .n32282(n32282), .n13576(n13576), .prev_select_adj_291(prev_select_adj_675), 
            .n32165(n32165), .n34065(n34065), .n34064(n34064), .n29977(n29977), 
            .n224({n224_adj_1021}), .n32(n32_adj_572), .n28053(n28053), 
            .read_value({read_value_adj_1017}), .n7062(n7033[3]), .n21184(n21184), 
            .n21176(n21176), .n29860(n29860), .\div_factor_reg[3] (div_factor_reg_adj_1015[3]), 
            .\databus[8] (databus[8]), .\databus[12] (databus[12]), .\databus[14] (databus[14]), 
            .int_step(int_step), .n22(n22_adj_571), .n32145(n32145), .n32153(n32153), 
            .n8585(n8584[7]), .n29983(n29983), .n14555(n14555)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(610[25] 623[45])
    ClockDivider_U10 pwm_clk_div (.n34065(n34065), .n7822(n7822), .n30615(n30615), 
            .n28233(n28233), .n30621(n30621), .n28222(n28222), .n30619(n30619), 
            .n28231(n28231), .debug_c_c(debug_c_c), .n241(n241), .n30482(n30482), 
            .n13605(n13605), .GND_net(battery_voltage[15]), .n32135(n32135), 
            .n30472(n30472), .n13974(n13974), .n30613(n30613), .n28234(n28234), 
            .n30623(n30623), .n28140(n28140), .n30617(n30617), .n28232(n28232), 
            .n30470(n30470), .n13975(n13975), .n30465(n30465), .n13976(n13976), 
            .n30463(n30463), .n13977(n13977), .n30474(n30474), .n32134(n32134)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(540[15] 543[41])
    \ArmPeripheral(axis_haddr=8'b010000)  arm_y (.debug_c_c(debug_c_c), .n34070(n34070), 
            .n34069(n34069), .\register_addr[0] (register_addr[0]), .VCC_net(VCC_net), 
            .GND_net(battery_voltage[15]), .Stepper_Y_nFault_c(Stepper_Y_nFault_c), 
            .n34066(n34066), .\read_size[0] (read_size_adj_980[0]), .n2776(n2776), 
            .n29713(n29713), .Stepper_Y_M0_c_0(Stepper_Y_M0_c_0), .n13899(n13899), 
            .n579(n571[0]), .prev_step_clk(prev_step_clk_adj_640), .step_clk(step_clk_adj_639), 
            .n13885(n13885), .prev_select(prev_select_adj_675), .n32163(n32163), 
            .read_value({read_value_adj_979}), .Stepper_Y_Step_c(Stepper_Y_Step_c), 
            .n32140(n32140), .n34067(n34067), .databus({databus}), .n34071(n34071), 
            .n608(n580_adj_998[4]), .\control_reg[7] (control_reg_adj_976[7]), 
            .n13576(n13576), .Stepper_Y_En_c(Stepper_Y_En_c), .Stepper_Y_Dir_c(Stepper_Y_Dir_c), 
            .Stepper_Y_M2_c_2(Stepper_Y_M2_c_2), .Stepper_Y_M1_c_1(Stepper_Y_M1_c_1), 
            .n4034(n4034), .\read_size[2] (read_size_adj_980[2]), .n28426(n28426), 
            .n34068(n34068), .\register_addr[1] (register_addr[1]), .limit_c_1(limit_c_1), 
            .n34065(n34065), .n32(n32), .n22(n22), .n32144(n32144), 
            .n8576(n8575[7]), .n28049(n28049)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(595[25] 608[45])
    LUT4 i20_2_lut_rep_320_3_lut_4_lut (.A(select[4]), .B(n32199), .C(rw), 
         .D(n32261), .Z(n32141)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i20_2_lut_rep_320_3_lut_4_lut.init = 16'h2000;
    CCU2D add_31_21 (.A0(timeout_count[19]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[20]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27040), 
          .COUT(n27041), .S0(n658[19]), .S1(n658[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_21.INIT0 = 16'h5aaa;
    defparam add_31_21.INIT1 = 16'h5aaa;
    defparam add_31_21.INJECT1_0 = "NO";
    defparam add_31_21.INJECT1_1 = "NO";
    RCPeripheral rc_receiver (.n2(n2_adj_681), .databus({databus}), .\register_addr[0] (register_addr[0]), 
            .\read_value[25] (read_value_adj_1055[25]), .n8(n8_adj_679), 
            .n32141(n32141), .n2_adj_58(n2_adj_725), .databus_out({databus_out}), 
            .n34064(n34064), .read_value({read_value_adj_979}), .\read_value[9]_adj_60 (read_value_adj_1100[9]), 
            .n52(n52_adj_676), .n32164(n32164), .\select[7] (select[7]), 
            .n176(n176), .n2_adj_61(n2_adj_569), .n2_adj_62(n2_adj_584), 
            .\read_value[11]_adj_63 (read_value_adj_1055[11]), .n8_adj_64(n8_adj_683), 
            .read_value_adj_287({read_value}), .read_value_adj_288({read_value_adj_967}), 
            .n46(n46), .n52_adj_129(n52), .\read_value[21]_adj_130 (read_value_adj_1055[21]), 
            .n8_adj_131(n8_adj_682), .n2_adj_132(n2_adj_677), .\read_value[20]_adj_133 (read_value_adj_1055[20]), 
            .n8_adj_134(n8_adj_934), .\read_value[11]_adj_135 (read_value_adj_1100[11]), 
            .rw(rw), .\read_value[20]_adj_136 (read_value_adj_1100[20]), 
            .read_size({read_size}), .\select[1] (select[1]), .n32284(n32284), 
            .\sendcount[1] (sendcount[1]), .n12746(n12746), .n2_adj_137(n2_adj_933), 
            .\read_value[19]_adj_138 (read_value_adj_1055[19]), .n8_adj_139(n8_adj_932), 
            .\register_addr[1] (register_addr[1]), .\read_value[19]_adj_140 (read_value_adj_1100[19]), 
            .n2_adj_141(n2_adj_809), .\read_value[10]_adj_142 (read_value_adj_1055[10]), 
            .n8_adj_143(n8_adj_846), .n3(n3_adj_882), .n2_adj_144(n2_adj_806), 
            .\read_value[18]_adj_145 (read_value_adj_1055[18]), .n8_adj_146(n8_adj_636), 
            .read_value_adj_289({read_value_adj_960}), .n64(n64), .n19559(n19559), 
            .read_value_adj_290({read_value_adj_1116}), .n2_adj_163(n2_adj_925), 
            .\read_value[18]_adj_164 (read_value_adj_1100[18]), .\read_value[3]_adj_165 (read_value_adj_1100[3]), 
            .\read_value[3]_adj_166 (read_value_adj_1092[3]), .n32161(n32161), 
            .n2_adj_167(n2_adj_845), .\read_value[8]_adj_168 (read_value_adj_1055[8]), 
            .n8_adj_169(n8_adj_680), .n3_adj_170(n3_adj_924), .n2_adj_171(n2_adj_580), 
            .\read_value[17]_adj_172 (read_value_adj_1055[17]), .n8_adj_173(n8_adj_902), 
            .\read_value[28]_adj_174 (read_value_adj_1055[28]), .n8_adj_175(n8_adj_907), 
            .\read_value[10]_adj_176 (read_value_adj_1100[10]), .\read_value[17]_adj_177 (read_value_adj_1100[17]), 
            .\register_addr[2] (register_addr[2]), .\register_addr[5] (register_addr[5]), 
            .n2_adj_178(n2_adj_586), .\read_value[16]_adj_179 (read_value_adj_1055[16]), 
            .n8_adj_180(n8_adj_582), .\read_value[16]_adj_181 (read_value_adj_1100[16]), 
            .\read_value[13]_adj_182 (read_value_adj_1100[13]), .\read_value[8]_adj_183 (read_value_adj_1100[8]), 
            .n2_adj_184(n2_adj_901), .\read_value[15]_adj_185 (read_value_adj_1055[15]), 
            .n8_adj_186(n8_adj_578), .\read_value[15]_adj_187 (read_value_adj_1100[15]), 
            .n32282(n32282), .\read_size[2]_adj_188 (read_size_adj_980[2]), 
            .\register_addr[4] (register_addr[4]), .\read_size[2]_adj_189 (read_size_adj_968[2]), 
            .n2_adj_190(n2_adj_929), .\read_value[2]_adj_191 (read_value_adj_1100[2]), 
            .\read_value[2]_adj_192 (read_value_adj_1092[2]), .\read_size[2]_adj_193 (read_size_adj_1018[2]), 
            .\read_size[2]_adj_194 (read_size_adj_1056[2]), .n2_adj_195(n2_adj_897), 
            .\read_value[14]_adj_196 (read_value_adj_1055[14]), .n8_adj_197(n8_adj_896), 
            .n3_adj_198(n3_adj_928), .n10(n10_adj_930), .\read_value[12]_adj_199 (read_value_adj_1055[12]), 
            .n8_adj_200(n8_adj_570), .\read_value[1]_adj_201 (read_value_adj_1092[1]), 
            .n3_adj_202(n3_adj_931), .\read_value[1]_adj_203 (read_value_adj_1055[1]), 
            .\read_value[14]_adj_204 (read_value_adj_1100[14]), .n2_adj_205(n2_adj_635), 
            .\read_value[9]_adj_206 (read_value_adj_1055[9]), .n8_adj_207(n8_adj_727), 
            .n2_adj_208(n2_adj_724), .\read_value[13]_adj_209 (read_value_adj_1055[13]), 
            .n8_adj_210(n8_adj_573), .\read_value[25]_adj_211 (read_value_adj_1100[25]), 
            .\read_value[28]_adj_212 (read_value_adj_1100[28]), .n2_adj_213(n2_adj_903), 
            .\read_value[27]_adj_214 (read_value_adj_1055[27]), .n8_adj_215(n8_adj_585), 
            .\read_value[27]_adj_216 (read_value_adj_1100[27]), .\read_value[21]_adj_217 (read_value_adj_1100[21]), 
            .n2_adj_218(n2_adj_919), .\read_value[6]_adj_219 (read_value_adj_1100[6]), 
            .\read_value[6]_adj_220 (read_value_adj_1092[6]), .n2_adj_221(n2_adj_637), 
            .n32185(n32185), .\read_value[24]_adj_222 (read_value_adj_1055[24]), 
            .n8_adj_223(n8_adj_684), .n13(n13_adj_895), .\read_size[0]_adj_224 (read_size_adj_1018[0]), 
            .n9(n9_adj_923), .n32215(n32215), .n18(n18), .\read_size[0]_adj_225 (read_size_adj_1093[0]), 
            .\read_size[0]_adj_226 (read_size_adj_961[0]), .n32182(n32182), 
            .\select[2] (select[2]), .n14(n14_adj_894), .\read_size[0]_adj_227 (read_size_adj_1056[0]), 
            .n5(n5), .n32155(n32155), .\read_size[0]_adj_228 (read_size_adj_1117[0]), 
            .\read_size[0]_adj_229 (read_size_adj_968[0]), .\select[5] (select[5]), 
            .n32203(n32203), .n32178(n32178), .\read_size[2]_adj_230 (read_size_adj_1101[2]), 
            .\reg_size[2] (reg_size[2]), .n3_adj_231(n3_adj_900), .\read_size[2]_adj_232 (read_size_adj_1093[2]), 
            .n32251(n32251), .n2_adj_233(n2_adj_597), .\read_value[26]_adj_234 (read_value_adj_1055[26]), 
            .n8_adj_235(n8_adj_921), .\read_value[26]_adj_236 (read_value_adj_1100[26]), 
            .\read_value[24]_adj_237 (read_value_adj_1100[24]), .\read_value[12]_adj_238 (read_value_adj_1100[12]), 
            .n2_adj_239(n2_adj_927), .\read_value[0]_adj_240 (read_value_adj_1100[0]), 
            .\read_value[0]_adj_241 (read_value_adj_1092[0]), .n3_adj_242(n3_adj_926), 
            .n2_adj_243(n2_adj_598), .\read_value[31]_adj_244 (read_value_adj_1055[31]), 
            .n8_adj_245(n8_adj_918), .\read_value[31]_adj_246 (read_value_adj_1100[31]), 
            .n2_adj_247(n2_adj_807), .n2_adj_248(n2_adj_583), .n2_adj_249(n2_adj_883), 
            .n29920(n29920), .n2_adj_250(n2_adj_579), .\read_value[30]_adj_251 (read_value_adj_1055[30]), 
            .n8_adj_252(n8_adj_568), .\read_value[30]_adj_253 (read_value_adj_1100[30]), 
            .\read_value[7]_adj_254 (read_value_adj_1100[7]), .\read_value[7]_adj_255 (read_value_adj_1092[7]), 
            .n2_adj_256(n2_adj_904), .\read_value[29]_adj_257 (read_value_adj_1055[29]), 
            .n8_adj_258(n8_adj_922), .\read_value[29]_adj_259 (read_value_adj_1100[29]), 
            .\read_value[4]_adj_260 (read_value_adj_1100[4]), .\read_value[4]_adj_261 (read_value_adj_1092[4]), 
            .n2_adj_262(n2_adj_905), .\read_value[5]_adj_263 (read_value_adj_1100[5]), 
            .\read_value[5]_adj_264 (read_value_adj_1092[5]), .\read_value[23]_adj_265 (read_value_adj_1055[23]), 
            .n8_adj_266(n8_adj_678), .\read_value[23]_adj_267 (read_value_adj_1100[23]), 
            .n3_adj_268(n3), .n3_adj_269(n3_adj_906), .n2_adj_270(n2_adj_808), 
            .\read_value[22]_adj_271 (read_value_adj_1055[22]), .n8_adj_272(n8), 
            .\read_value[22]_adj_273 (read_value_adj_1100[22]), .n2_adj_274(n2), 
            .\count[6] (count_adj_1267[6]), .\count[5] (count_adj_1267[5]), 
            .n29947(n29947), .n5_adj_275(n5_adj_917), .GND_net(battery_voltage[15]), 
            .n30260(n30260), .\count[8] (count_adj_1267[8]), .\count[9] (count_adj_1267[9]), 
            .n30482(n30482), .n32135(n32135), .n30304(n30304), .n32302(n32302), 
            .\count[4] (count_adj_1267[4]), .n32245(n32245), .n32301(n32301), 
            .n28333(n28333), .debug_c_c(debug_c_c), .rc_ch8_c(rc_ch8_c), 
            .n32256(n32256), .\count[1] (count_adj_1267[1]), .\count[2] (count_adj_1267[2]), 
            .n32257(n32257), .\count[3] (count_adj_1267[3]), .n32218(n32218), 
            .n32258(n32258), .n13605(n13605), .\count[0] (count_adj_1267[0]), 
            .n30001(n30001), .n29948(n29948), .n28141(n28141), .n28234(n28234), 
            .n32129(n32129), .n32134(n32134), .n30474(n30474), .rc_ch7_c(rc_ch7_c), 
            .n30623(n30623), .n28140(n28140), .n32283(n32283), .n28331(n28331), 
            .n32317(n32317), .n13974(n13974), .rc_ch4_c(rc_ch4_c), .n28133(n28133), 
            .n30472(n30472), .n28233(n28233), .n32221(n32221), .\count[9]_adj_276 (count_adj_1228[9]), 
            .n32264(n32264), .n28330(n28330), .n5_adj_277(n5_adj_912), 
            .\count[5]_adj_278 (count_adj_1228[5]), .n5_adj_279(n5_adj_599), 
            .\count[6]_adj_280 (count_adj_1228[6]), .n32267(n32267), .\count[8]_adj_281 (count_adj_1228[8]), 
            .n13975(n13975), .rc_ch3_c(rc_ch3_c), .n28132(n28132), .n28222(n28222), 
            .n32127(n32127), .n30470(n30470), .n30302(n30302), .n28232(n28232), 
            .n32125(n32125), .n32294(n32294), .\count[9]_adj_282 (count_adj_1215[9]), 
            .\count[8]_adj_283 (count_adj_1215[8]), .\count[5]_adj_284 (count_adj_1215[5]), 
            .\count[6]_adj_285 (count_adj_1215[6]), .rc_ch2_c(rc_ch2_c), 
            .n13976(n13976), .n5_adj_286(n5_adj_920), .n32293(n32293), 
            .n41(n41), .n28329(n28329), .n32296(n32296), .n28144(n28144), 
            .n30308(n30308), .n30465(n30465), .n13977(n13977), .n30463(n30463), 
            .n32274(n32274), .n28328(n28328), .n32308(n32308), .rc_ch1_c(rc_ch1_c), 
            .n28231(n28231), .n28129(n28129)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(708[15] 720[41])
    CCU2D add_31_19 (.A0(timeout_count[17]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[18]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27039), 
          .COUT(n27040), .S0(n658[17]), .S1(n658[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_19.INIT0 = 16'h5aaa;
    defparam add_31_19.INIT1 = 16'h5aaa;
    defparam add_31_19.INJECT1_0 = "NO";
    defparam add_31_19.INJECT1_1 = "NO";
    CCU2D add_31_17 (.A0(timeout_count[15]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[16]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27038), 
          .COUT(n27039), .S0(n658[15]), .S1(n658[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_17.INIT0 = 16'h5aaa;
    defparam add_31_17.INIT1 = 16'h5aaa;
    defparam add_31_17.INJECT1_0 = "NO";
    defparam add_31_17.INJECT1_1 = "NO";
    LUT4 i14756_3_lut (.A(Stepper_A_En_c), .B(div_factor_reg_adj_1053[6]), 
         .C(register_addr[1]), .Z(n21445)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i14756_3_lut.init = 16'hcaca;
    SabertoothSerialPeripheral motor_serial (.debug_c_c(debug_c_c), .n13545(n13545), 
            .n282(n281[15]), .n32147(n32147), .n34066(n34066), .\databus[6] (databus[6]), 
            .n34070(n34070), .\databus[5] (databus[5]), .\databus[4] (databus[4]), 
            .n34067(n34067), .\databus[3] (databus[3]), .\databus[2] (databus[2]), 
            .\databus[1] (databus[1]), .\databus[0] (databus[0]), .\register[0] ({\register[0]_adj_959 [7], 
            Open_0, Open_1, Open_2, Open_3, Open_4, Open_5, Open_6}), 
            .n13560(n13560), .n32146(n32146), .\read_size[0] (read_size_adj_961[0]), 
            .n2760(n2760), .n21718(n21718), .n34068(n34068), .prev_select(prev_select_adj_596), 
            .\select[2] (select[2]), .\register_addr[0] (register_addr[0]), 
            .n32285(n32285), .read_value({read_value_adj_960}), .n9482(n9482), 
            .GND_net(battery_voltage[15]), .n34065(n34065), .n8447(n8447), 
            .n32227(n32227), .state({state_adj_1287}), .n29194(n29194), 
            .n11013(n11013), .n34071(n34071), .n29883(n29883), .n107(n107)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(530[29] 538[56])
    \ClockDividerP_SP(factor=120000)  clk_100Hz_divider (.debug_c_0(debug_c_0), 
            .debug_c_c(debug_c_c), .n34070(n34070), .n34065(n34065), .GND_net(battery_voltage[15])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(643[29] 645[61])
    GlobalControlPeripheral global_control (.read_value({read_value}), .debug_c_c(debug_c_c), 
            .n14419(n14419), .n9478(n9478), .n34068(n34068), .read_size({read_size}), 
            .n302(n302), .prev_select(prev_select), .\select[1] (select[1]), 
            .n28365(n28365), .n13412(n13412), .n34065(n34065), .n34066(n34066), 
            .n34070(n34070), .n34071(n34071), .\register_addr[0] (register_addr[0]), 
            .\register_addr[1] (register_addr[1]), .timeout_pause(timeout_pause), 
            .n32285(n32285), .\register[0][7] (\register[0]_adj_959 [7]), 
            .n32227(n32227), .signal_light_c(signal_light_c), .rw(rw), 
            .n46(n46), .n16516(n16516), .n30075(n30075), .n16515(n16515), 
            .n32158(n32158), .n32200(n32200), .xbee_pause_c(xbee_pause_c), 
            .GND_net(battery_voltage[15]), .n34067(n34067), .\databus[1] (databus[1]), 
            .n30270(n30270), .n34069(n34069)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(514[45] 525[74])
    LUT4 i23217_4_lut (.A(n32274), .B(n32308), .C(n28328), .D(n28129), 
         .Z(n30619)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;
    defparam i23217_4_lut.init = 16'h5455;
    LUT4 i14753_3_lut (.A(control_reg_adj_1052[3]), .B(div_factor_reg_adj_1053[3]), 
         .C(register_addr[1]), .Z(n21442)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i14753_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_493 (.A(register_addr[1]), .B(n9496), .Z(n29758)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_2_lut_adj_493.init = 16'h2222;
    LUT4 i1_4_lut_adj_494 (.A(div_factor_reg_adj_1053[9]), .B(n29758), .C(steps_reg_adj_1054[9]), 
         .D(register_addr[0]), .Z(n29759)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_4_lut_adj_494.init = 16'hc088;
    LUT4 i14488_3_lut (.A(Stepper_Z_Dir_c), .B(div_factor_reg_adj_1015[5]), 
         .C(register_addr[1]), .Z(n21182)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i14488_3_lut.init = 16'hcaca;
    EncoderPeripheral_U11 left_encoder (.read_value({read_value_adj_1092}), 
            .debug_c_c(debug_c_c), .n14271(n14271), .n32160(n32160), .\read_size[0] (read_size_adj_1093[0]), 
            .n302(n302), .\quadA_delayed[1] (quadA_delayed_adj_1199[1]), 
            .qreset(qreset), .n6(n6), .\quadB_delayed[1] (quadB_delayed_adj_1200[1]), 
            .n13588(n13588), .n34065(n34065), .debug_c_0(debug_c_0), .prev_select(prev_select_adj_844), 
            .n32182(n32182), .n32232(n32232), .n32235(n32235), .n32278(n32278), 
            .n9482(n9482), .\register_addr[0] (register_addr[0]), .encoder_li_c(encoder_li_c), 
            .encoder_lb_c(encoder_lb_c), .encoder_la_c(encoder_la_c), .\read_size[2] (read_size_adj_1093[2]), 
            .n32158(n32158), .VCC_net(VCC_net), .GND_net(battery_voltage[15])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(671[20] 681[47])
    LUT4 i23211_4_lut (.A(n5_adj_917), .B(n32301), .C(n28333), .D(n28141), 
         .Z(n30613)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;
    defparam i23211_4_lut.init = 16'h5455;
    LUT4 i1_4_lut_adj_495 (.A(count_adj_1228[8]), .B(n32267), .C(count_adj_1228[5]), 
         .D(n32221), .Z(n44_adj_726)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_adj_495.init = 16'heaaa;
    LUT4 i23160_3_lut (.A(count_adj_1228[8]), .B(count_adj_1228[6]), .C(n5_adj_599), 
         .Z(n30324)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i23160_3_lut.init = 16'h0101;
    VLO i1 (.Z(battery_voltage[15]));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i23087_4_lut_4_lut (.A(n32213), .B(n4), .C(n5774), .D(n1414[14]), 
         .Z(n13567)) /* synthesis lut_function=(!((B (C+!(D))+!B !(D))+!A)) */ ;
    defparam i23087_4_lut_4_lut.init = 16'h2a00;
    LUT4 i14480_3_lut (.A(Stepper_Z_En_c), .B(div_factor_reg_adj_1015[6]), 
         .C(register_addr[1]), .Z(n21174)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i14480_3_lut.init = 16'hcaca;
    LUT4 i8_2_lut (.A(timeout_count[1]), .B(timeout_count[4]), .Z(n30_adj_899)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i18_4_lut (.A(timeout_count[6]), .B(n36), .C(n26), .D(timeout_count[2]), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i14477_3_lut (.A(control_reg_adj_1014[3]), .B(div_factor_reg_adj_1015[3]), 
         .C(register_addr[1]), .Z(n21171)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i14477_3_lut.init = 16'hcaca;
    PFUMX i14766 (.BLUT(n21453), .ALUT(n14), .C0(register_addr[0]), .Z(n21455));
    CCU2D add_31_15 (.A0(timeout_count[13]), .B0(battery_voltage[15]), .C0(battery_voltage[15]), 
          .D0(battery_voltage[15]), .A1(timeout_count[14]), .B1(battery_voltage[15]), 
          .C1(battery_voltage[15]), .D1(battery_voltage[15]), .CIN(n27037), 
          .COUT(n27038), .S0(n658[13]), .S1(n658[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(482[24:41])
    defparam add_31_15.INIT0 = 16'h5aaa;
    defparam add_31_15.INIT1 = 16'h5aaa;
    defparam add_31_15.INJECT1_0 = "NO";
    defparam add_31_15.INJECT1_1 = "NO";
    PFUMX i14758 (.BLUT(n21445), .ALUT(n13), .C0(register_addr[0]), .Z(n21447));
    \ProtocolInterface(baud_div=12)  protocol_interface (.register_addr({register_addr}), 
            .debug_c_c(debug_c_c), .n13118(n13118), .n29983(n29983), .databus({databus}), 
            .n224({n224_adj_1059}), .n3862({n3862}), .debug_c_7(debug_c_7), 
            .n32213(n32213), .n32261(n32261), .n32235(n32235), .n32315(n32315), 
            .n29712(n29712), .\select[5] (select[5]), .rw(rw), .n19559(n19559), 
            .n32152(n32152), .n34064(n34064), .n13567(n13567), .databus_out({databus_out}), 
            .\sendcount[1] (sendcount[1]), .n32153(n32153), .n224_adj_56({n224_adj_1021}), 
            .n3948({n3948}), .n32172(n32172), .n32278(n32278), .n34065(n34065), 
            .n13560(n13560), .\select[7] (select[7]), .\select[4] (select[4]), 
            .\select[3] (select[3]), .\select[2] (select[2]), .\select[1] (select[1]), 
            .n1432(n1414[14]), .n13545(n13545), .prev_select(prev_select_adj_596), 
            .n2760(n2760), .n32279(n32279), .n29750(n29750), .n32154(n32154), 
            .n13885(n13885), .n21718(n21718), .n32282(n32282), .n32233(n32233), 
            .n32202(n32202), .n32231(n32231), .n32137(n32137), .n32253(n32253), 
            .n112(n112), .n30075(n30075), .debug_c_5(debug_c_5), .n32251(n32251), 
            .n52(n52), .prev_select_adj_41(prev_select_adj_634), .n32181(n32181), 
            .n32305(n32305), .n32182(n32182), .n29713(n29713), .n32178(n32178), 
            .n5774(n5774), .n32314(n32314), .n28302(n28302), .n32316(n32316), 
            .n32252(n32252), .n13576(n13576), .n13899(n13899), .n32165(n32165), 
            .n13769(n13769), .\control_reg[7] (control_reg_adj_1014[7]), 
            .n8585(n8584[7]), .n32168(n32168), .prev_select_adj_42(prev_select_adj_675), 
            .n32163(n32163), .n32140(n32140), .n29977(n29977), .n4034(n4034), 
            .n64(n64), .\control_reg[7]_adj_43 (control_reg_adj_1052[7]), 
            .n8594(n8593[7]), .\control_reg[7]_adj_44 (control_reg[7]), 
            .n1(n1), .n12746(n12746), .n13(n13_adj_895), .n18(n18), 
            .n14(n14_adj_894), .n32155(n32155), .\reg_size[2] (reg_size[2]), 
            .n32284(n32284), .n28062(n28062), .n32285(n32285), .n34(n34), 
            .n28053(n28053), .n32(n32_adj_572), .debug_c_2(debug_c_2), 
            .debug_c_3(debug_c_3), .debug_c_4(debug_c_4), .\steps_reg[5] (steps_reg_adj_1054[5]), 
            .n14_adj_45(n14), .n28049(n28049), .\control_reg[7]_adj_46 (control_reg_adj_976[7]), 
            .n32_adj_47(n32), .\steps_reg[6] (steps_reg_adj_1054[6]), .n13_adj_48(n13), 
            .\steps_reg[3] (steps_reg_adj_1054[3]), .n12(n12), .n4(n4), 
            .n28061(n28061), .n32_adj_49(n32_adj_574), .\steps_reg[5]_adj_50 (steps_reg_adj_1016[5]), 
            .n14_adj_51(n14_adj_577), .\steps_reg[6]_adj_52 (steps_reg_adj_1016[6]), 
            .n13_adj_53(n13_adj_576), .n32234(n32234), .n13412(n13412), 
            .\steps_reg[3]_adj_54 (steps_reg_adj_1016[3]), .n12_adj_55(n12_adj_581), 
            .n8576(n8575[7]), .\reset_count[14] (reset_count[14]), .\reset_count[13] (reset_count[13]), 
            .\reset_count[12] (reset_count[12]), .n29954(n29954), .uart_tx_c(uart_tx_c), 
            .GND_net(battery_voltage[15]), .uart_rx_c(uart_rx_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(493[26] 503[57])
    LUT4 i1_4_lut_adj_496 (.A(count_adj_1267[8]), .B(n32258), .C(count_adj_1267[5]), 
         .D(n32218), .Z(n44)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_adj_496.init = 16'heaaa;
    PFUMX i14755 (.BLUT(n21442), .ALUT(n12), .C0(register_addr[0]), .Z(n7347[3]));
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_497 (.A(n34065), .B(prev_select_adj_675), 
         .C(n32168), .D(n32305), .Z(n2776)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_497.init = 16'h1000;
    LUT4 i15306_2_lut_2_lut (.A(n34065), .B(databus[0]), .Z(n571[0])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i15306_2_lut_2_lut.init = 16'h4444;
    LUT4 i23172_3_lut (.A(count_adj_1267[8]), .B(count_adj_1267[6]), .C(n30260), 
         .Z(n30330)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i23172_3_lut.init = 16'h0101;
    LUT4 i12_4_lut (.A(timeout_count[14]), .B(timeout_count[11]), .C(timeout_count[30]), 
         .D(timeout_count[13]), .Z(n34_adj_898)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(timeout_count[29]), .B(timeout_count[26]), .C(timeout_count[7]), 
         .D(timeout_count[3]), .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(timeout_count[0]), .B(timeout_count[27]), .Z(n26)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(485[7:35])
    defparam i4_2_lut.init = 16'heeee;
    PFUMX i14490 (.BLUT(n21182), .ALUT(n14_adj_577), .C0(register_addr[0]), 
          .Z(n21184));
    \ArmPeripheral(axis_haddr=8'b0)  arm_x (.databus({databus}), .debug_c_c(debug_c_c), 
            .n34069(n34069), .n608(n580_adj_998[4]), .n610(n580_adj_1036[2]), 
            .\control_reg[7] (control_reg[7]), .n32149(n32149), .Stepper_X_En_c(Stepper_X_En_c), 
            .Stepper_X_Dir_c(Stepper_X_Dir_c), .n13511(n13511), .Stepper_X_M2_c_2(Stepper_X_M2_c_2), 
            .Stepper_X_M1_c_1(Stepper_X_M1_c_1), .\read_size[2] (read_size_adj_968[2]), 
            .n2769(n2769), .n21617(n21617), .n34067(n34067), .n34068(n34068), 
            .n34071(n34071), .\read_size[0] (read_size_adj_968[0]), .n21718(n21718), 
            .n34066(n34066), .Stepper_X_M0_c_0(Stepper_X_M0_c_0), .n579(n571[0]), 
            .prev_step_clk(prev_step_clk), .step_clk(step_clk), .prev_select(prev_select_adj_634), 
            .n32203(n32203), .read_value({read_value_adj_967}), .n9485(n9485), 
            .Stepper_X_Step_c(Stepper_X_Step_c), .\register_addr[1] (register_addr[1]), 
            .\register_addr[0] (register_addr[0]), .rw(rw), .n32181(n32181), 
            .n32233(n32233), .n29750(n29750), .n32279(n32279), .n13118(n13118), 
            .n32231(n32231), .n32235(n32235), .n32232(n32232), .n22529(n22529), 
            .n14812(n14812), .n32282(n32282), .n32314(n32314), .n32315(n32315), 
            .n30020(n30020), .n32305(n32305), .n28426(n28426), .n32261(n32261), 
            .n30019(n30019), .n32187(n32187), .limit_c_0(limit_c_0), .n32159(n32159), 
            .n34065(n34065), .n14419(n14419), .n9478(n9478), .n1(n1), 
            .n34(n34), .n28062(n28062), .VCC_net(VCC_net), .GND_net(battery_voltage[15]), 
            .Stepper_X_nFault_c(Stepper_X_nFault_c), .n24(n24), .n32142(n32142)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(580[25] 593[45])
    CCU2D reset_count_2657_2658_add_4_15 (.A0(reset_count[13]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[14]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27397), .S0(n66_adj_1469[13]), .S1(n66_adj_1469[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658_add_4_15.INIT0 = 16'hfaaa;
    defparam reset_count_2657_2658_add_4_15.INIT1 = 16'hfaaa;
    defparam reset_count_2657_2658_add_4_15.INJECT1_0 = "NO";
    defparam reset_count_2657_2658_add_4_15.INJECT1_1 = "NO";
    CCU2D reset_count_2657_2658_add_4_13 (.A0(reset_count[11]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[12]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27396), .COUT(n27397), .S0(n66_adj_1469[11]), .S1(n66_adj_1469[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658_add_4_13.INIT0 = 16'hfaaa;
    defparam reset_count_2657_2658_add_4_13.INIT1 = 16'hfaaa;
    defparam reset_count_2657_2658_add_4_13.INJECT1_0 = "NO";
    defparam reset_count_2657_2658_add_4_13.INJECT1_1 = "NO";
    EncoderPeripheral right_encoder (.\read_size[0] (read_size_adj_1101[0]), 
            .debug_c_c(debug_c_c), .n178(n178), .n32157(n32157), .n32202(n32202), 
            .read_value({read_value_adj_1100}), .prev_select(prev_select_adj_881), 
            .n32178(n32178), .\register_addr[0] (register_addr[0]), .n32235(n32235), 
            .n32232(n32232), .prev_select_adj_8(prev_select), .n30270(n30270), 
            .n32315(n32315), .n29983(n29983), .n32138(n32138), .n29977(n29977), 
            .n9(n9), .\read_size[2] (read_size_adj_1101[2]), .\register_addr[1] (register_addr[1]), 
            .n32282(n32282), .n32166(n32166), .n32279(n32279), .n32204(n32204), 
            .n32181(n32181), .rw(rw), .n32149(n32149), .n34065(n34065), 
            .n32159(n32159), .n13511(n13511), .encoder_ra_c(encoder_ra_c), 
            .encoder_rb_c(encoder_rb_c), .encoder_ri_c(encoder_ri_c), .n14493(n14493), 
            .n14419(n14419), .n32231(n32231), .n16516(n16516), .n16515(n16515), 
            .n6(n6), .n13588(n13588), .qreset(qreset), .VCC_net(VCC_net), 
            .GND_net(battery_voltage[15]), .\quadB_delayed[1] (quadB_delayed_adj_1200[1]), 
            .\quadA_delayed[1] (quadA_delayed_adj_1199[1])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(682[20] 692[47])
    \ArmPeripheral(axis_haddr=8'b0110000)  arm_a (.Stepper_A_M0_c_0(Stepper_A_M0_c_0), 
            .\register_addr[0] (register_addr[0]), .debug_c_c(debug_c_c), 
            .n34066(n34066), .n3862({n3862}), .VCC_net(VCC_net), .GND_net(battery_voltage[15]), 
            .Stepper_A_nFault_c(Stepper_A_nFault_c), .\read_size[0] (read_size_adj_1056[0]), 
            .n14114(n14114), .n29712(n29712), .n14493(n14493), .n579(n571[0]), 
            .n14555(n14555), .prev_select(prev_select_adj_773), .n32155(n32155), 
            .\read_size[2] (read_size_adj_1056[2]), .n30019(n30019), .n34068(n34068), 
            .Stepper_A_M1_c_1(Stepper_A_M1_c_1), .n34069(n34069), .\steps_reg[9] (steps_reg_adj_1054[9]), 
            .\steps_reg[6] (steps_reg_adj_1054[6]), .\steps_reg[5] (steps_reg_adj_1054[5]), 
            .\steps_reg[3] (steps_reg_adj_1054[3]), .n34065(n34065), .prev_step_clk(prev_step_clk), 
            .n34(n34), .step_clk(step_clk), .n32142(n32142), .n24(n24), 
            .n32(n32_adj_574), .n32_adj_1(n32), .prev_step_clk_adj_2(prev_step_clk_adj_640), 
            .step_clk_adj_3(step_clk_adj_639), .n32144(n32144), .limit_c_3(limit_c_3), 
            .n22(n22), .n32_adj_4(n32_adj_572), .prev_step_clk_adj_5(prev_step_clk_adj_687), 
            .step_clk_adj_6(step_clk_adj_686), .n32145(n32145), .n22_adj_7(n22_adj_571), 
            .n224({n224_adj_1059}), .\register_addr[1] (register_addr[1]), 
            .n32138(n32138), .n34071(n34071), .\databus[1] (databus[1]), 
            .Stepper_A_M2_c_2(Stepper_A_M2_c_2), .n610(n580_adj_1036[2]), 
            .\control_reg[3] (control_reg_adj_1052[3]), .\databus[3] (databus[3]), 
            .n608(n580_adj_998[4]), .Stepper_A_Dir_c(Stepper_A_Dir_c), .\databus[5] (databus[5]), 
            .Stepper_A_En_c(Stepper_A_En_c), .\databus[6] (databus[6]), 
            .\control_reg[7] (control_reg_adj_1052[7]), .\databus[7] (databus[7]), 
            .\div_factor_reg[5] (div_factor_reg_adj_1053[5]), .n32137(n32137), 
            .\div_factor_reg[6] (div_factor_reg_adj_1053[6]), .\div_factor_reg[9] (div_factor_reg_adj_1053[9]), 
            .\databus[9] (databus[9]), .\databus[10] (databus[10]), .\databus[11] (databus[11]), 
            .\databus[13] (databus[13]), .n32216(n32216), .\databus[22] (databus[22]), 
            .\databus[23] (databus[23]), .\databus[24] (databus[24]), .\databus[25] (databus[25]), 
            .\databus[26] (databus[26]), .\databus[27] (databus[27]), .\databus[28] (databus[28]), 
            .\databus[29] (databus[29]), .\databus[30] (databus[30]), .\databus[31] (databus[31]), 
            .\databus[21] (databus[21]), .\databus[20] (databus[20]), .\databus[19] (databus[19]), 
            .\databus[18] (databus[18]), .\databus[17] (databus[17]), .\databus[16] (databus[16]), 
            .\databus[15] (databus[15]), .\databus[14] (databus[14]), .\databus[12] (databus[12]), 
            .\databus[8] (databus[8]), .\div_factor_reg[3] (div_factor_reg_adj_1053[3]), 
            .int_step(int_step_adj_738), .read_value({read_value_adj_1055}), 
            .n9496(n9496), .n7376(n7347[3]), .n21455(n21455), .n21447(n21447), 
            .n29759(n29759), .n8594(n8593[7]), .n29758(n29758), .n28061(n28061)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(625[25] 638[45])
    LUT4 i15001_2_lut_2_lut (.A(n34065), .B(n7822), .Z(n241)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i15001_2_lut_2_lut.init = 16'h4444;
    CCU2D reset_count_2657_2658_add_4_11 (.A0(reset_count[9]), .B0(battery_voltage[15]), 
          .C0(battery_voltage[15]), .D0(battery_voltage[15]), .A1(reset_count[10]), 
          .B1(battery_voltage[15]), .C1(battery_voltage[15]), .D1(battery_voltage[15]), 
          .CIN(n27395), .COUT(n27396), .S0(n66_adj_1469[9]), .S1(n66_adj_1469[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[20:35])
    defparam reset_count_2657_2658_add_4_11.INIT0 = 16'hfaaa;
    defparam reset_count_2657_2658_add_4_11.INIT1 = 16'hfaaa;
    defparam reset_count_2657_2658_add_4_11.INJECT1_0 = "NO";
    defparam reset_count_2657_2658_add_4_11.INJECT1_1 = "NO";
    PFUMX i14482 (.BLUT(n21174), .ALUT(n13_adj_576), .C0(register_addr[0]), 
          .Z(n21176));
    PFUMX i14479 (.BLUT(n21171), .ALUT(n12_adj_581), .C0(register_addr[0]), 
          .Z(n7033[3]));
    
endmodule
//
// Verilog Description of module ExpansionGPIO
//

module ExpansionGPIO (read_value, debug_c_c, n32162, n13598, n34066, 
            \databus[0] , \read_size[0] , n22529, prev_select, \select[5] , 
            n10948, n10947, expansion1_c_9, n14812, expansion2_c_10, 
            expansion3_c_11, expansion5_c, n32187, n32204, \register_addr[0] , 
            expansion4_out, n32315, n32279, n32235, n302, n32158, 
            rw, n32172, \register_addr[1] , n32282, n21617, n32278, 
            n32146, n32147, n32306, n32216, \databus[1] , \databus[2] , 
            \databus[3] , \databus[4] , \databus[5] , \databus[6] , 
            \databus[7] , n11961, n16718, n32232, \register_addr[3] , 
            n29920, \register_addr[2] , n176, n32185, n112, n28365) /* synthesis syn_module_defined=1 */ ;
    output [7:0]read_value;
    input debug_c_c;
    input n32162;
    input n13598;
    input n34066;
    input \databus[0] ;
    output \read_size[0] ;
    input n22529;
    output prev_select;
    input \select[5] ;
    output n10948;
    output n10947;
    output expansion1_c_9;
    input n14812;
    output expansion2_c_10;
    output expansion3_c_11;
    input expansion5_c;
    input n32187;
    input n32204;
    input \register_addr[0] ;
    input expansion4_out;
    input n32315;
    input n32279;
    input n32235;
    output n302;
    output n32158;
    input rw;
    output n32172;
    input \register_addr[1] ;
    input n32282;
    output n21617;
    input n32278;
    output n32146;
    output n32147;
    input n32306;
    input n32216;
    input \databus[1] ;
    input \databus[2] ;
    input \databus[3] ;
    input \databus[4] ;
    input \databus[5] ;
    input \databus[6] ;
    input \databus[7] ;
    input n11961;
    input n16718;
    input n32232;
    input \register_addr[3] ;
    input n29920;
    input \register_addr[2] ;
    output n176;
    output n32185;
    input n112;
    output n28365;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [7:0]n7577;
    wire [7:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(17[12:20])
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(17[12:20])
    
    wire n30262;
    wire [7:0]n7602;
    
    wire n15085;
    
    FD1P3AX read_value_i0_i4 (.D(n7577[4]), .SP(n32162), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i4.GSR = "ENABLED";
    FD1P3IX register_0___i1 (.D(\databus[0] ), .SP(n13598), .CD(n34066), 
            .CK(debug_c_c), .Q(\register[0] [0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i1.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n22529), .SP(n32162), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1S3AX prev_select_145 (.D(\select[5] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam prev_select_145.GSR = "ENABLED";
    LUT4 Select_4204_i3_4_lut (.A(\register[1] [4]), .B(\register[1] [5]), 
         .C(\register[0] [4]), .D(\register[0] [5]), .Z(n10948)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam Select_4204_i3_4_lut.init = 16'heca0;
    LUT4 i23151_2_lut (.A(\register[0] [5]), .B(\register[0] [4]), .Z(n10947)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i23151_2_lut.init = 16'h1111;
    LUT4 mux_2016_i2_4_lut (.A(expansion1_c_9), .B(\register[0] [1]), .C(n14812), 
         .D(n30262), .Z(n7577[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2016_i2_4_lut.init = 16'ha0ac;
    LUT4 mux_2016_i3_4_lut (.A(expansion2_c_10), .B(\register[0] [2]), .C(n14812), 
         .D(n30262), .Z(n7577[2])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2016_i3_4_lut.init = 16'ha0ac;
    LUT4 mux_2016_i4_4_lut (.A(expansion3_c_11), .B(\register[0] [3]), .C(n14812), 
         .D(n30262), .Z(n7577[3])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2016_i4_4_lut.init = 16'ha0ac;
    LUT4 mux_2016_i6_4_lut (.A(expansion5_c), .B(n7602[5]), .C(n32187), 
         .D(n32204), .Z(n7577[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2016_i6_4_lut.init = 16'h0aca;
    LUT4 mux_2017_Mux_5_i1_3_lut (.A(\register[0] [5]), .B(\register[1] [5]), 
         .C(\register_addr[0] ), .Z(n7602[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2017_Mux_5_i1_3_lut.init = 16'hcaca;
    LUT4 mux_2016_i5_4_lut (.A(expansion4_out), .B(n7602[4]), .C(n32187), 
         .D(n32204), .Z(n7577[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2016_i5_4_lut.init = 16'h0aca;
    LUT4 mux_2017_Mux_4_i1_3_lut (.A(\register[0] [4]), .B(\register[1] [4]), 
         .C(\register_addr[0] ), .Z(n7602[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2017_Mux_4_i1_3_lut.init = 16'hcaca;
    LUT4 equal_138_i16_1_lut_2_lut_2_lut_3_lut_4_lut (.A(n32315), .B(n32279), 
         .C(n32235), .D(\register_addr[0] ), .Z(n302)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(116[11:28])
    defparam equal_138_i16_1_lut_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 equal_138_i15_2_lut_rep_337_2_lut_3_lut_4_lut (.A(n32315), .B(n32279), 
         .C(n32235), .D(\register_addr[0] ), .Z(n32158)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(116[11:28])
    defparam equal_138_i15_2_lut_rep_337_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i15003_2_lut_rep_351_3_lut_4_lut (.A(n32315), .B(n32279), .C(rw), 
         .D(n32235), .Z(n32172)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(116[11:28])
    defparam i15003_2_lut_rep_351_3_lut_4_lut.init = 16'hfffe;
    LUT4 i23055_2_lut_2_lut_3_lut_4_lut (.A(n32315), .B(n32279), .C(\register_addr[1] ), 
         .D(n32282), .Z(n21617)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(116[11:28])
    defparam i23055_2_lut_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i22759_2_lut_3_lut_4_lut (.A(n32315), .B(n32279), .C(\register_addr[0] ), 
         .D(n32235), .Z(n30262)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(116[11:28])
    defparam i22759_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_325_3_lut_4_lut (.A(rw), .B(n32204), .C(\register_addr[0] ), 
         .D(n32278), .Z(n32146)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_325_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_326_3_lut_4_lut (.A(rw), .B(n32204), .C(\register_addr[0] ), 
         .D(n32278), .Z(n32147)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_326_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut (.A(rw), .B(n32204), .C(\register_addr[0] ), 
         .D(n32306), .Z(n15085)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 mux_2017_Mux_7_i1_3_lut (.A(\register[0] [7]), .B(\register[1] [7]), 
         .C(\register_addr[0] ), .Z(n7602[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2017_Mux_7_i1_3_lut.init = 16'hcaca;
    LUT4 mux_2017_Mux_6_i1_3_lut (.A(\register[0] [6]), .B(\register[1] [6]), 
         .C(\register_addr[0] ), .Z(n7602[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2017_Mux_6_i1_3_lut.init = 16'hcaca;
    FD1P3IX register_0___i2 (.D(\databus[1] ), .SP(n13598), .CD(n32216), 
            .CK(debug_c_c), .Q(\register[0] [1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i2.GSR = "ENABLED";
    FD1P3IX register_0___i3 (.D(\databus[2] ), .SP(n13598), .CD(n32216), 
            .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i3.GSR = "ENABLED";
    FD1P3IX register_0___i4 (.D(\databus[3] ), .SP(n13598), .CD(n32216), 
            .CK(debug_c_c), .Q(\register[0] [3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i4.GSR = "ENABLED";
    FD1P3IX register_0___i5 (.D(\databus[4] ), .SP(n13598), .CD(n32216), 
            .CK(debug_c_c), .Q(\register[0] [4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i5.GSR = "ENABLED";
    FD1P3IX register_0___i6 (.D(\databus[5] ), .SP(n13598), .CD(n32216), 
            .CK(debug_c_c), .Q(\register[0] [5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i6.GSR = "ENABLED";
    FD1P3IX register_0___i7 (.D(\databus[6] ), .SP(n13598), .CD(n32216), 
            .CK(debug_c_c), .Q(\register[0] [6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i7.GSR = "ENABLED";
    FD1P3IX register_0___i8 (.D(\databus[7] ), .SP(n13598), .CD(n32216), 
            .CK(debug_c_c), .Q(\register[0] [7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i8.GSR = "ENABLED";
    FD1P3IX register_0___i9 (.D(\databus[0] ), .SP(n15085), .CD(n32216), 
            .CK(debug_c_c), .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i9.GSR = "ENABLED";
    FD1P3IX register_0___i10 (.D(\databus[1] ), .SP(n15085), .CD(n32216), 
            .CK(debug_c_c), .Q(expansion1_c_9)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i10.GSR = "ENABLED";
    FD1P3IX register_0___i11 (.D(\databus[2] ), .SP(n11961), .CD(n32216), 
            .CK(debug_c_c), .Q(expansion2_c_10)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i11.GSR = "ENABLED";
    FD1P3IX register_0___i12 (.D(\databus[3] ), .SP(n11961), .CD(n32216), 
            .CK(debug_c_c), .Q(expansion3_c_11)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i12.GSR = "ENABLED";
    FD1P3IX register_0___i13 (.D(\databus[4] ), .SP(n11961), .CD(n32216), 
            .CK(debug_c_c), .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i13.GSR = "ENABLED";
    FD1P3IX register_0___i14 (.D(\databus[5] ), .SP(n11961), .CD(n32216), 
            .CK(debug_c_c), .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i14.GSR = "ENABLED";
    FD1P3IX register_0___i15 (.D(\databus[6] ), .SP(n11961), .CD(n32216), 
            .CK(debug_c_c), .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i15.GSR = "ENABLED";
    FD1P3IX register_0___i16 (.D(\databus[7] ), .SP(n11961), .CD(n32216), 
            .CK(debug_c_c), .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam register_0___i16.GSR = "ENABLED";
    FD1P3AX read_value_i0_i1 (.D(n7577[1]), .SP(n32162), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i1.GSR = "ENABLED";
    FD1P3AX read_value_i0_i2 (.D(n7577[2]), .SP(n32162), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i2.GSR = "ENABLED";
    FD1P3AX read_value_i0_i3 (.D(n7577[3]), .SP(n32162), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i3.GSR = "ENABLED";
    FD1P3AX read_value_i0_i5 (.D(n7577[5]), .SP(n32162), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i5.GSR = "ENABLED";
    FD1P3IX read_value_i0_i7 (.D(n7602[7]), .SP(n32162), .CD(n16718), 
            .CK(debug_c_c), .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i7.GSR = "ENABLED";
    FD1P3IX read_value_i0_i6 (.D(n7602[6]), .SP(n32162), .CD(n16718), 
            .CK(debug_c_c), .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i6.GSR = "ENABLED";
    LUT4 i15936_1_lut_3_lut_4_lut (.A(n32232), .B(\register_addr[3] ), .C(n29920), 
         .D(\register_addr[2] ), .Z(n176)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;
    defparam i15936_1_lut_3_lut_4_lut.init = 16'h0111;
    LUT4 i1_3_lut_rep_364_4_lut (.A(n32232), .B(\register_addr[3] ), .C(n29920), 
         .D(\register_addr[2] ), .Z(n32185)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_3_lut_rep_364_4_lut.init = 16'hfeee;
    FD1P3IX read_value_i0_i0 (.D(n7602[0]), .SP(n32162), .CD(n16718), 
            .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=38, LSE_LLINE=694, LSE_RLINE=705 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(34[9] 77[6])
    defparam read_value_i0_i0.GSR = "ENABLED";
    LUT4 mux_2017_Mux_0_i1_3_lut (.A(\register[0] [0]), .B(\register[1] [0]), 
         .C(\register_addr[0] ), .Z(n7602[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/expansion.v(45[7] 66[14])
    defparam mux_2017_Mux_0_i1_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(n32232), .B(\register_addr[3] ), .C(\register_addr[2] ), 
         .D(n112), .Z(n28365)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hffef;
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0100000) 
//

module \ArmPeripheral(axis_haddr=8'b0100000)  (limit_c_2, Stepper_Z_M0_c_0, 
            register_addr, debug_c_c, VCC_net, GND_net, Stepper_Z_nFault_c, 
            n34066, n3948, \read_size[0] , n13476, n28302, n579, 
            prev_step_clk, step_clk, n13769, prev_select, n32215, 
            n34067, \databus[31] , \databus[30] , \databus[29] , \databus[28] , 
            \databus[27] , \databus[26] , \databus[25] , \databus[24] , 
            \databus[23] , \databus[22] , \databus[21] , \databus[20] , 
            \databus[19] , \databus[18] , \databus[17] , \databus[16] , 
            \databus[15] , n34068, \databus[13] , \databus[11] , \databus[10] , 
            \div_factor_reg[9] , \databus[9] , \databus[7] , \div_factor_reg[6] , 
            \databus[6] , \div_factor_reg[5] , \databus[5] , n608, n610, 
            \control_reg[7] , Stepper_Z_En_c, Stepper_Z_Dir_c, \control_reg[3] , 
            \databus[3] , Stepper_Z_M2_c_2, Stepper_Z_M1_c_1, \databus[1] , 
            \read_size[2] , n30020, n34070, \steps_reg[9] , \steps_reg[6] , 
            n34071, \steps_reg[5] , \steps_reg[3] , n32315, n29750, 
            n32232, n32234, n32316, n32200, n32205, \select[4] , 
            n32251, n32253, rw, n32189, n32252, n32199, n32166, 
            n32314, n9, n32282, n13576, prev_select_adj_291, n32165, 
            n34065, n34064, n29977, n224, n32, n28053, read_value, 
            n7062, n21184, n21176, n29860, \div_factor_reg[3] , \databus[8] , 
            \databus[12] , \databus[14] , int_step, n22, n32145, n32153, 
            n8585, n29983, n14555) /* synthesis syn_module_defined=1 */ ;
    input limit_c_2;
    output Stepper_Z_M0_c_0;
    input [7:0]register_addr;
    input debug_c_c;
    input VCC_net;
    input GND_net;
    input Stepper_Z_nFault_c;
    input n34066;
    input [31:0]n3948;
    output \read_size[0] ;
    input n13476;
    input n28302;
    input n579;
    output prev_step_clk;
    output step_clk;
    input n13769;
    output prev_select;
    input n32215;
    input n34067;
    input \databus[31] ;
    input \databus[30] ;
    input \databus[29] ;
    input \databus[28] ;
    input \databus[27] ;
    input \databus[26] ;
    input \databus[25] ;
    input \databus[24] ;
    input \databus[23] ;
    input \databus[22] ;
    input \databus[21] ;
    input \databus[20] ;
    input \databus[19] ;
    input \databus[18] ;
    input \databus[17] ;
    input \databus[16] ;
    input \databus[15] ;
    input n34068;
    input \databus[13] ;
    input \databus[11] ;
    input \databus[10] ;
    output \div_factor_reg[9] ;
    input \databus[9] ;
    input \databus[7] ;
    output \div_factor_reg[6] ;
    input \databus[6] ;
    output \div_factor_reg[5] ;
    input \databus[5] ;
    input n608;
    input n610;
    output \control_reg[7] ;
    output Stepper_Z_En_c;
    output Stepper_Z_Dir_c;
    output \control_reg[3] ;
    input \databus[3] ;
    output Stepper_Z_M2_c_2;
    output Stepper_Z_M1_c_1;
    input \databus[1] ;
    output \read_size[2] ;
    input n30020;
    input n34070;
    output \steps_reg[9] ;
    output \steps_reg[6] ;
    input n34071;
    output \steps_reg[5] ;
    output \steps_reg[3] ;
    output n32315;
    output n29750;
    output n32232;
    output n32234;
    input n32316;
    output n32200;
    output n32205;
    input \select[4] ;
    output n32251;
    output n32253;
    input rw;
    input n32189;
    input n32252;
    output n32199;
    input n32166;
    input n32314;
    input n9;
    input n32282;
    output n13576;
    input prev_select_adj_291;
    input n32165;
    input n34065;
    input n34064;
    output n29977;
    output [31:0]n224;
    input n32;
    output n28053;
    output [31:0]read_value;
    input n7062;
    input n21184;
    input n21176;
    input n29860;
    output \div_factor_reg[3] ;
    input \databus[8] ;
    input \databus[12] ;
    input \databus[14] ;
    output int_step;
    input n22;
    input n32145;
    output n32153;
    input n8585;
    input n29983;
    output n14555;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n182, limit_latched, n30351;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire n30352, fault_latched, n13823, prev_limit_latched, n32151, 
        n32139, n11176;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [7:0]n8584;
    
    wire n30402, n30403, n30404;
    wire [31:0]n6997;
    
    wire n30198, n30353, n27462, n27461, n27460, n30363, n30364, 
        n27459, n30365, n27458, n27457, n27456, n27455, n27454, 
        n27453, n27452, n27451, n27450, n27449, n27448, n27447, 
        n49, n62, n58, n50;
    wire [31:0]n7033;
    
    wire n29861, n29862, n29863, n29864, n29865, n29866, n29867, 
        n29868, n29869, n29870, n29871, n29872, n29857, n29859, 
        n29873, n29874, n29875, n29876, n29877, n29878, n29879, 
        n29880, n41, n60, n54, n42, n52, n38, n29858, n56, 
        n46;
    
    LUT4 i118_1_lut (.A(limit_c_2), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i22848_3_lut (.A(Stepper_Z_M0_c_0), .B(limit_latched), .C(register_addr[0]), 
         .Z(n30351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22848_3_lut.init = 16'hcaca;
    LUT4 i22849_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(register_addr[0]), 
         .Z(n30352)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22849_3_lut.init = 16'hcaca;
    IFS1P3DX fault_latched_178 (.D(Stepper_Z_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3948[0]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n28302), .SP(n13476), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n13823), .CK(debug_c_c), .Q(Stepper_Z_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n13769), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n32215), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(\databus[31] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(\databus[30] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(\databus[29] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(\databus[28] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(\databus[27] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(\databus[26] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(\databus[25] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(\databus[24] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(\databus[23] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(\databus[22] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(\databus[21] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(\databus[20] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(\databus[19] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(\databus[18] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(\databus[17] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(\databus[16] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(\databus[15] ), .SP(n32151), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(\databus[13] ), .SP(n32151), .PD(n34068), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(\databus[11] ), .SP(n32151), .PD(n34068), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(\databus[10] ), .SP(n32151), .PD(n34068), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(\databus[9] ), .SP(n32151), .PD(n34068), 
            .CK(debug_c_c), .Q(\div_factor_reg[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(\databus[7] ), .SP(n32151), .PD(n34068), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(\databus[6] ), .SP(n32151), .PD(n34068), 
            .CK(debug_c_c), .Q(\div_factor_reg[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(\databus[5] ), .SP(n32151), .PD(n34068), 
            .CK(debug_c_c), .Q(\div_factor_reg[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n13769), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n13769), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(\databus[7] ), .SP(n32139), .CD(n11176), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(\databus[6] ), .SP(n32139), .PD(n34068), 
            .CK(debug_c_c), .Q(Stepper_Z_En_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(\databus[5] ), .SP(n32139), .PD(n34068), 
            .CK(debug_c_c), .Q(Stepper_Z_Dir_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n13823), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(\databus[3] ), .SP(n32139), .PD(n34068), 
            .CK(debug_c_c), .Q(\control_reg[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n13823), .CK(debug_c_c), .Q(Stepper_Z_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(\databus[1] ), .SP(n32139), .PD(n34068), 
            .CK(debug_c_c), .Q(Stepper_Z_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    LUT4 i15259_2_lut (.A(control_reg[4]), .B(register_addr[0]), .Z(n8584[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15259_2_lut.init = 16'h2222;
    FD1P3AX read_size__i2 (.D(n30020), .SP(n13476), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3948[31]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3948[30]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3948[29]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3948[28]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3948[27]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3948[26]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3948[25]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3948[24]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3948[23]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3948[22]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3948[21]), .CK(debug_c_c), .CD(n34067), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3948[20]), .CK(debug_c_c), .CD(n34067), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3948[19]), .CK(debug_c_c), .CD(n34067), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3948[18]), .CK(debug_c_c), .CD(n34067), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3948[17]), .CK(debug_c_c), .CD(n34067), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3948[16]), .CK(debug_c_c), .CD(n34067), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3948[15]), .CK(debug_c_c), .CD(n34067), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3948[14]), .CK(debug_c_c), .CD(n34067), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3948[13]), .CK(debug_c_c), .CD(n34067), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3948[12]), .CK(debug_c_c), .CD(n34067), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3948[11]), .CK(debug_c_c), .CD(n34067), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3948[10]), .CK(debug_c_c), .CD(n34070), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3948[9]), .CK(debug_c_c), .CD(n34070), 
            .Q(\steps_reg[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3948[8]), .CK(debug_c_c), .CD(n34070), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3948[7]), .CK(debug_c_c), .CD(n34070), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3948[6]), .CK(debug_c_c), .CD(n34071), 
            .Q(\steps_reg[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3948[5]), .CK(debug_c_c), .CD(n34070), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3948[4]), .CK(debug_c_c), .CD(n34070), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3948[3]), .CK(debug_c_c), .CD(n34070), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3948[2]), .CK(debug_c_c), .CD(n34071), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3948[1]), .CK(debug_c_c), .CD(n34070), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    PFUMX i22901 (.BLUT(n30402), .ALUT(n30403), .C0(register_addr[0]), 
          .Z(n30404));
    LUT4 i1_2_lut_rep_494 (.A(register_addr[6]), .B(register_addr[7]), .Z(n32315)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_494.init = 16'heeee;
    LUT4 i1_3_lut_4_lut (.A(register_addr[6]), .B(register_addr[7]), .C(register_addr[0]), 
         .D(register_addr[1]), .Z(n29750)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_411_3_lut_4_lut (.A(register_addr[6]), .B(register_addr[7]), 
         .C(register_addr[4]), .D(register_addr[5]), .Z(n32232)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_411_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_413_3_lut (.A(register_addr[6]), .B(register_addr[7]), 
         .C(register_addr[5]), .Z(n32234)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_413_3_lut.init = 16'hfefe;
    LUT4 mux_1964_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(register_addr[0]), 
         .Z(n6997[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1964_i5_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_379_3_lut_4_lut (.A(register_addr[6]), .B(register_addr[7]), 
         .C(n32316), .D(register_addr[5]), .Z(n32200)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_379_3_lut_4_lut.init = 16'hfffe;
    LUT4 i4374_2_lut_rep_384_3_lut_4_lut (.A(register_addr[6]), .B(register_addr[7]), 
         .C(register_addr[4]), .D(register_addr[5]), .Z(n32205)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i4374_2_lut_rep_384_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_430_3_lut (.A(register_addr[6]), .B(register_addr[7]), 
         .C(\select[4] ), .Z(n32251)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_430_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_rep_432_3_lut (.A(register_addr[6]), .B(register_addr[7]), 
         .C(register_addr[3]), .Z(n32253)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_432_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_rep_330_4_lut (.A(rw), .B(n32189), .C(n29750), .D(n32252), 
         .Z(n32151)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i2_3_lut_rep_330_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_rep_378_3_lut_4_lut (.A(register_addr[6]), .B(register_addr[7]), 
         .C(register_addr[2]), .D(register_addr[3]), .Z(n32199)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_378_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_318_3_lut_4_lut (.A(rw), .B(n32189), .C(n32166), 
         .D(n32314), .Z(n32139)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i1_2_lut_rep_318_3_lut_4_lut.init = 16'h0004;
    LUT4 i5_4_lut (.A(n9), .B(n30198), .C(n32282), .D(\select[4] ), 
         .Z(n13576)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(83[9:13])
    defparam i5_4_lut.init = 16'h0200;
    LUT4 i22699_2_lut (.A(register_addr[5]), .B(prev_select_adj_291), .Z(n30198)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22699_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32165), .B(n32314), .C(n34065), .D(n32166), 
         .Z(n13823)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(83[9:13])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf0f2;
    LUT4 i1_2_lut (.A(n34064), .B(register_addr[4]), .Z(n29977)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(83[9:13])
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i4460_3_lut (.A(prev_limit_latched), .B(n34065), .C(limit_latched), 
         .Z(n11176)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i4460_3_lut.init = 16'hdcdc;
    LUT4 mux_1964_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(register_addr[0]), 
         .Z(n6997[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1964_i8_3_lut.init = 16'hcaca;
    PFUMX i22850 (.BLUT(n30351), .ALUT(n30352), .C0(register_addr[1]), 
          .Z(n30353));
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27462), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27461), .COUT(n27462), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27460), .COUT(n27461), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    LUT4 i22860_3_lut (.A(Stepper_Z_M1_c_1), .B(fault_latched), .C(register_addr[0]), 
         .Z(n30363)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22860_3_lut.init = 16'hcaca;
    LUT4 i22861_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(register_addr[0]), 
         .Z(n30364)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22861_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27459), .COUT(n27460), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    PFUMX i22862 (.BLUT(n30363), .ALUT(n30364), .C0(register_addr[1]), 
          .Z(n30365));
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27458), .COUT(n27459), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27457), .COUT(n27458), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27456), .COUT(n27457), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27455), .COUT(n27456), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27454), .COUT(n27455), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27453), .COUT(n27454), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27452), .COUT(n27453), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(\steps_reg[9] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27451), .COUT(n27452), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27450), .COUT(n27451), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27449), .COUT(n27450), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27448), .COUT(n27449), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27447), .COUT(n27448), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n27447), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i22899_3_lut (.A(Stepper_Z_M2_c_2), .B(div_factor_reg[2]), .C(register_addr[1]), 
         .Z(n30402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22899_3_lut.init = 16'hcaca;
    LUT4 i22900_3_lut (.A(n32), .B(steps_reg[2]), .C(register_addr[1]), 
         .Z(n30403)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22900_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n28053)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[0]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    FD1P3IX read_value__i1 (.D(n30365), .SP(n13476), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30404), .SP(n13476), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n7062), .SP(n13476), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n7033[4]), .SP(n13476), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n21184), .SP(n13476), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n21176), .SP(n13476), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n7033[7]), .SP(n13476), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29861), .SP(n13476), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29860), .SP(n13476), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29862), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29863), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29864), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29865), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29866), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29867), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29868), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29869), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29870), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n29871), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29872), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29857), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(\databus[1] ), .SP(n13769), .CD(n34068), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29859), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29873), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(\databus[3] ), .SP(n13769), .CD(n34068), 
            .CK(debug_c_c), .Q(\div_factor_reg[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29874), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(\databus[8] ), .SP(n13769), .CD(n34068), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n29875), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(\databus[12] ), .SP(n13769), .CD(n34068), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(\databus[14] ), .SP(n13769), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n29876), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n29877), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n29878), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n29879), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n29880), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52), .C(n38), .D(steps_reg[18]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    FD1P3AX read_value__i31 (.D(n29858), .SP(n13476), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX int_step_182 (.D(n32145), .SP(n22), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n30353), .SP(n13476), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=610, LSE_RLINE=623 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i9_2_lut (.A(steps_reg[7]), .B(\steps_reg[5] ), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[26]), .B(n56), .C(n46), .D(steps_reg[29]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[25]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[10]), .B(steps_reg[22]), .C(steps_reg[20]), 
         .D(\steps_reg[6] ), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(\steps_reg[9] ), .B(\steps_reg[3] ), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[28]), .C(steps_reg[13]), 
         .D(steps_reg[30]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[2]), .B(steps_reg[8]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i1_4_lut (.A(div_factor_reg[8]), .B(register_addr[1]), .C(steps_reg[8]), 
         .D(register_addr[0]), .Z(n29861)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_460 (.A(div_factor_reg[10]), .B(register_addr[1]), 
         .C(steps_reg[10]), .D(register_addr[0]), .Z(n29862)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_460.init = 16'hc088;
    LUT4 i1_4_lut_adj_461 (.A(div_factor_reg[11]), .B(register_addr[1]), 
         .C(steps_reg[11]), .D(register_addr[0]), .Z(n29863)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_461.init = 16'hc088;
    LUT4 i1_4_lut_adj_462 (.A(div_factor_reg[12]), .B(register_addr[1]), 
         .C(steps_reg[12]), .D(register_addr[0]), .Z(n29864)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_462.init = 16'hc088;
    LUT4 i1_4_lut_adj_463 (.A(div_factor_reg[13]), .B(register_addr[1]), 
         .C(steps_reg[13]), .D(register_addr[0]), .Z(n29865)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_463.init = 16'hc088;
    LUT4 i1_4_lut_adj_464 (.A(div_factor_reg[14]), .B(register_addr[1]), 
         .C(steps_reg[14]), .D(register_addr[0]), .Z(n29866)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_464.init = 16'hc088;
    LUT4 i1_4_lut_adj_465 (.A(div_factor_reg[15]), .B(register_addr[1]), 
         .C(steps_reg[15]), .D(register_addr[0]), .Z(n29867)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_465.init = 16'hc088;
    LUT4 i1_4_lut_adj_466 (.A(div_factor_reg[16]), .B(register_addr[1]), 
         .C(steps_reg[16]), .D(register_addr[0]), .Z(n29868)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_466.init = 16'hc088;
    LUT4 i1_4_lut_adj_467 (.A(div_factor_reg[17]), .B(register_addr[1]), 
         .C(steps_reg[17]), .D(register_addr[0]), .Z(n29869)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_467.init = 16'hc088;
    LUT4 i1_4_lut_adj_468 (.A(div_factor_reg[18]), .B(register_addr[1]), 
         .C(steps_reg[18]), .D(register_addr[0]), .Z(n29870)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_468.init = 16'hc088;
    LUT4 i1_4_lut_adj_469 (.A(div_factor_reg[19]), .B(register_addr[1]), 
         .C(steps_reg[19]), .D(register_addr[0]), .Z(n29871)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_469.init = 16'hc088;
    LUT4 i1_4_lut_adj_470 (.A(div_factor_reg[20]), .B(register_addr[1]), 
         .C(steps_reg[20]), .D(register_addr[0]), .Z(n29872)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_470.init = 16'hc088;
    LUT4 i1_4_lut_adj_471 (.A(div_factor_reg[21]), .B(register_addr[1]), 
         .C(steps_reg[21]), .D(register_addr[0]), .Z(n29857)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_471.init = 16'hc088;
    LUT4 i1_4_lut_adj_472 (.A(div_factor_reg[22]), .B(register_addr[1]), 
         .C(steps_reg[22]), .D(register_addr[0]), .Z(n29859)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_472.init = 16'hc088;
    LUT4 i1_4_lut_adj_473 (.A(div_factor_reg[23]), .B(register_addr[1]), 
         .C(steps_reg[23]), .D(register_addr[0]), .Z(n29873)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_473.init = 16'hc088;
    LUT4 i1_4_lut_adj_474 (.A(div_factor_reg[24]), .B(register_addr[1]), 
         .C(steps_reg[24]), .D(register_addr[0]), .Z(n29874)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_474.init = 16'hc088;
    LUT4 i1_4_lut_adj_475 (.A(div_factor_reg[25]), .B(register_addr[1]), 
         .C(steps_reg[25]), .D(register_addr[0]), .Z(n29875)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_475.init = 16'hc088;
    LUT4 i1_4_lut_adj_476 (.A(div_factor_reg[26]), .B(register_addr[1]), 
         .C(steps_reg[26]), .D(register_addr[0]), .Z(n29876)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_476.init = 16'hc088;
    LUT4 i1_4_lut_adj_477 (.A(div_factor_reg[27]), .B(register_addr[1]), 
         .C(steps_reg[27]), .D(register_addr[0]), .Z(n29877)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_477.init = 16'hc088;
    LUT4 i1_4_lut_adj_478 (.A(div_factor_reg[28]), .B(register_addr[1]), 
         .C(steps_reg[28]), .D(register_addr[0]), .Z(n29878)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_478.init = 16'hc088;
    LUT4 i1_4_lut_adj_479 (.A(div_factor_reg[29]), .B(register_addr[1]), 
         .C(steps_reg[29]), .D(register_addr[0]), .Z(n29879)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_479.init = 16'hc088;
    LUT4 i1_4_lut_adj_480 (.A(div_factor_reg[30]), .B(register_addr[1]), 
         .C(steps_reg[30]), .D(register_addr[0]), .Z(n29880)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_480.init = 16'hc088;
    LUT4 i1_4_lut_adj_481 (.A(div_factor_reg[31]), .B(register_addr[1]), 
         .C(steps_reg[31]), .D(register_addr[0]), .Z(n29858)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_481.init = 16'hc088;
    LUT4 i1_2_lut_rep_332_3_lut_4_lut (.A(n32215), .B(prev_select), .C(n32314), 
         .D(n34064), .Z(n32153)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i1_2_lut_rep_332_3_lut_4_lut.init = 16'h0002;
    PFUMX mux_1968_i5 (.BLUT(n8584[4]), .ALUT(n6997[4]), .C0(register_addr[1]), 
          .Z(n7033[4]));
    PFUMX mux_1968_i8 (.BLUT(n8585), .ALUT(n6997[7]), .C0(register_addr[1]), 
          .Z(n7033[7]));
    LUT4 i1_2_lut_4_lut (.A(n29983), .B(n32282), .C(n29750), .D(n34065), 
         .Z(n14555)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;
    defparam i1_2_lut_4_lut.init = 16'hff20;
    ClockDivider step_clk_gen (.GND_net(GND_net), .step_clk(step_clk), .debug_c_c(debug_c_c), 
            .n34070(n34070), .div_factor_reg({div_factor_reg[31:10], \div_factor_reg[9] , 
            div_factor_reg[8:7], \div_factor_reg[6] , \div_factor_reg[5] , 
            div_factor_reg[4], \div_factor_reg[3] , div_factor_reg[2:0]}), 
            .n34065(n34065)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider
//

module ClockDivider (GND_net, step_clk, debug_c_c, n34070, div_factor_reg, 
            n34065) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output step_clk;
    input debug_c_c;
    input n34070;
    input [31:0]div_factor_reg;
    input n34065;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27511;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    wire [31:0]n40;
    
    wire n27512, n27214;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    
    wire n8169, n27213, n27212, n27211, n27210, n27209, n32132;
    wire [31:0]n134;
    
    wire n16806, n27208, n27207, n27206, n27205, n27204, n27203, 
        n27202, n27201, n27200, n27199, n27198, n8204, n27197, 
        n27196, n27195, n27194, n27193, n27192, n27191, n27190, 
        n27189, n27188, n27582, n27187, n27186, n27185, n27184, 
        n27581, n27183, n27182, n8238, n27181, n27580, n27180, 
        n27179, n27178, n27177, n27176, n27579, n27175, n27174, 
        n27578, n27577, n27576, n27173, n27172, n27171, n27575, 
        n27574, n27170, n27169, n27168, n27573, n27572, n27571, 
        n27167, n27570, n27569, n27568, n27567, n27526, n27525, 
        n27524, n27523, n27522, n27521, n27520, n27519, n27518, 
        n27517, n27516, n27515, n27514, n27513;
    
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27511), .COUT(n27512), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27511), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2062_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27214), .S1(n8169));
    defparam sub_2062_add_2_33.INIT0 = 16'h5555;
    defparam sub_2062_add_2_33.INIT1 = 16'h0000;
    defparam sub_2062_add_2_33.INJECT1_0 = "NO";
    defparam sub_2062_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2062_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27213), .COUT(n27214));
    defparam sub_2062_add_2_31.INIT0 = 16'h5999;
    defparam sub_2062_add_2_31.INIT1 = 16'h5999;
    defparam sub_2062_add_2_31.INJECT1_0 = "NO";
    defparam sub_2062_add_2_31.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n8169), .CK(debug_c_c), .CD(n34070), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2062_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27212), .COUT(n27213));
    defparam sub_2062_add_2_29.INIT0 = 16'h5999;
    defparam sub_2062_add_2_29.INIT1 = 16'h5999;
    defparam sub_2062_add_2_29.INJECT1_0 = "NO";
    defparam sub_2062_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2062_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27211), .COUT(n27212));
    defparam sub_2062_add_2_27.INIT0 = 16'h5999;
    defparam sub_2062_add_2_27.INIT1 = 16'h5999;
    defparam sub_2062_add_2_27.INJECT1_0 = "NO";
    defparam sub_2062_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2062_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27210), .COUT(n27211));
    defparam sub_2062_add_2_25.INIT0 = 16'h5999;
    defparam sub_2062_add_2_25.INIT1 = 16'h5999;
    defparam sub_2062_add_2_25.INJECT1_0 = "NO";
    defparam sub_2062_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2062_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27209), .COUT(n27210));
    defparam sub_2062_add_2_23.INIT0 = 16'h5999;
    defparam sub_2062_add_2_23.INIT1 = 16'h5999;
    defparam sub_2062_add_2_23.INJECT1_0 = "NO";
    defparam sub_2062_add_2_23.INJECT1_1 = "NO";
    FD1S3IX count_2664__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i0.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    CCU2D sub_2062_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27208), .COUT(n27209));
    defparam sub_2062_add_2_21.INIT0 = 16'h5999;
    defparam sub_2062_add_2_21.INIT1 = 16'h5999;
    defparam sub_2062_add_2_21.INJECT1_0 = "NO";
    defparam sub_2062_add_2_21.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n32132), .PD(n16806), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_2062_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27207), .COUT(n27208));
    defparam sub_2062_add_2_19.INIT0 = 16'h5999;
    defparam sub_2062_add_2_19.INIT1 = 16'h5999;
    defparam sub_2062_add_2_19.INJECT1_0 = "NO";
    defparam sub_2062_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2062_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27206), .COUT(n27207));
    defparam sub_2062_add_2_17.INIT0 = 16'h5999;
    defparam sub_2062_add_2_17.INIT1 = 16'h5999;
    defparam sub_2062_add_2_17.INJECT1_0 = "NO";
    defparam sub_2062_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2062_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27205), .COUT(n27206));
    defparam sub_2062_add_2_15.INIT0 = 16'h5999;
    defparam sub_2062_add_2_15.INIT1 = 16'h5999;
    defparam sub_2062_add_2_15.INJECT1_0 = "NO";
    defparam sub_2062_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2062_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27204), .COUT(n27205));
    defparam sub_2062_add_2_13.INIT0 = 16'h5999;
    defparam sub_2062_add_2_13.INIT1 = 16'h5999;
    defparam sub_2062_add_2_13.INJECT1_0 = "NO";
    defparam sub_2062_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2062_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27203), .COUT(n27204));
    defparam sub_2062_add_2_11.INIT0 = 16'h5999;
    defparam sub_2062_add_2_11.INIT1 = 16'h5999;
    defparam sub_2062_add_2_11.INJECT1_0 = "NO";
    defparam sub_2062_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2062_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27202), .COUT(n27203));
    defparam sub_2062_add_2_9.INIT0 = 16'h5999;
    defparam sub_2062_add_2_9.INIT1 = 16'h5999;
    defparam sub_2062_add_2_9.INJECT1_0 = "NO";
    defparam sub_2062_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2062_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27201), .COUT(n27202));
    defparam sub_2062_add_2_7.INIT0 = 16'h5999;
    defparam sub_2062_add_2_7.INIT1 = 16'h5999;
    defparam sub_2062_add_2_7.INJECT1_0 = "NO";
    defparam sub_2062_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2062_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27200), .COUT(n27201));
    defparam sub_2062_add_2_5.INIT0 = 16'h5999;
    defparam sub_2062_add_2_5.INIT1 = 16'h5999;
    defparam sub_2062_add_2_5.INJECT1_0 = "NO";
    defparam sub_2062_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2062_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27199), .COUT(n27200));
    defparam sub_2062_add_2_3.INIT0 = 16'h5999;
    defparam sub_2062_add_2_3.INIT1 = 16'h5999;
    defparam sub_2062_add_2_3.INJECT1_0 = "NO";
    defparam sub_2062_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2062_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27199));
    defparam sub_2062_add_2_1.INIT0 = 16'h0000;
    defparam sub_2062_add_2_1.INIT1 = 16'h5999;
    defparam sub_2062_add_2_1.INJECT1_0 = "NO";
    defparam sub_2062_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27198), .S1(n8204));
    defparam sub_2064_add_2_33.INIT0 = 16'h5999;
    defparam sub_2064_add_2_33.INIT1 = 16'h0000;
    defparam sub_2064_add_2_33.INJECT1_0 = "NO";
    defparam sub_2064_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27197), .COUT(n27198));
    defparam sub_2064_add_2_31.INIT0 = 16'h5999;
    defparam sub_2064_add_2_31.INIT1 = 16'h5999;
    defparam sub_2064_add_2_31.INJECT1_0 = "NO";
    defparam sub_2064_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27196), .COUT(n27197));
    defparam sub_2064_add_2_29.INIT0 = 16'h5999;
    defparam sub_2064_add_2_29.INIT1 = 16'h5999;
    defparam sub_2064_add_2_29.INJECT1_0 = "NO";
    defparam sub_2064_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27195), .COUT(n27196));
    defparam sub_2064_add_2_27.INIT0 = 16'h5999;
    defparam sub_2064_add_2_27.INIT1 = 16'h5999;
    defparam sub_2064_add_2_27.INJECT1_0 = "NO";
    defparam sub_2064_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27194), .COUT(n27195));
    defparam sub_2064_add_2_25.INIT0 = 16'h5999;
    defparam sub_2064_add_2_25.INIT1 = 16'h5999;
    defparam sub_2064_add_2_25.INJECT1_0 = "NO";
    defparam sub_2064_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27193), .COUT(n27194));
    defparam sub_2064_add_2_23.INIT0 = 16'h5999;
    defparam sub_2064_add_2_23.INIT1 = 16'h5999;
    defparam sub_2064_add_2_23.INJECT1_0 = "NO";
    defparam sub_2064_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27192), .COUT(n27193));
    defparam sub_2064_add_2_21.INIT0 = 16'h5999;
    defparam sub_2064_add_2_21.INIT1 = 16'h5999;
    defparam sub_2064_add_2_21.INJECT1_0 = "NO";
    defparam sub_2064_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27191), .COUT(n27192));
    defparam sub_2064_add_2_19.INIT0 = 16'h5999;
    defparam sub_2064_add_2_19.INIT1 = 16'h5999;
    defparam sub_2064_add_2_19.INJECT1_0 = "NO";
    defparam sub_2064_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27190), .COUT(n27191));
    defparam sub_2064_add_2_17.INIT0 = 16'h5999;
    defparam sub_2064_add_2_17.INIT1 = 16'h5999;
    defparam sub_2064_add_2_17.INJECT1_0 = "NO";
    defparam sub_2064_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27189), .COUT(n27190));
    defparam sub_2064_add_2_15.INIT0 = 16'h5999;
    defparam sub_2064_add_2_15.INIT1 = 16'h5999;
    defparam sub_2064_add_2_15.INJECT1_0 = "NO";
    defparam sub_2064_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27188), .COUT(n27189));
    defparam sub_2064_add_2_13.INIT0 = 16'h5999;
    defparam sub_2064_add_2_13.INIT1 = 16'h5999;
    defparam sub_2064_add_2_13.INJECT1_0 = "NO";
    defparam sub_2064_add_2_13.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27582), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_33.INIT1 = 16'h0000;
    defparam count_2664_add_4_33.INJECT1_0 = "NO";
    defparam count_2664_add_4_33.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27187), .COUT(n27188));
    defparam sub_2064_add_2_11.INIT0 = 16'h5999;
    defparam sub_2064_add_2_11.INIT1 = 16'h5999;
    defparam sub_2064_add_2_11.INJECT1_0 = "NO";
    defparam sub_2064_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27186), .COUT(n27187));
    defparam sub_2064_add_2_9.INIT0 = 16'h5999;
    defparam sub_2064_add_2_9.INIT1 = 16'h5999;
    defparam sub_2064_add_2_9.INJECT1_0 = "NO";
    defparam sub_2064_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27185), .COUT(n27186));
    defparam sub_2064_add_2_7.INIT0 = 16'h5999;
    defparam sub_2064_add_2_7.INIT1 = 16'h5999;
    defparam sub_2064_add_2_7.INJECT1_0 = "NO";
    defparam sub_2064_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27184), .COUT(n27185));
    defparam sub_2064_add_2_5.INIT0 = 16'h5999;
    defparam sub_2064_add_2_5.INIT1 = 16'h5999;
    defparam sub_2064_add_2_5.INJECT1_0 = "NO";
    defparam sub_2064_add_2_5.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27581), .COUT(n27582), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2664_add_4_31.INJECT1_0 = "NO";
    defparam count_2664_add_4_31.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27183), .COUT(n27184));
    defparam sub_2064_add_2_3.INIT0 = 16'h5999;
    defparam sub_2064_add_2_3.INIT1 = 16'h5999;
    defparam sub_2064_add_2_3.INJECT1_0 = "NO";
    defparam sub_2064_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2064_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27183));
    defparam sub_2064_add_2_1.INIT0 = 16'h0000;
    defparam sub_2064_add_2_1.INIT1 = 16'h5999;
    defparam sub_2064_add_2_1.INJECT1_0 = "NO";
    defparam sub_2064_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27182), .S1(n8238));
    defparam sub_2065_add_2_33.INIT0 = 16'hf555;
    defparam sub_2065_add_2_33.INIT1 = 16'h0000;
    defparam sub_2065_add_2_33.INJECT1_0 = "NO";
    defparam sub_2065_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27181), .COUT(n27182));
    defparam sub_2065_add_2_31.INIT0 = 16'hf555;
    defparam sub_2065_add_2_31.INIT1 = 16'hf555;
    defparam sub_2065_add_2_31.INJECT1_0 = "NO";
    defparam sub_2065_add_2_31.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27580), .COUT(n27581), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2664_add_4_29.INJECT1_0 = "NO";
    defparam count_2664_add_4_29.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27180), .COUT(n27181));
    defparam sub_2065_add_2_29.INIT0 = 16'hf555;
    defparam sub_2065_add_2_29.INIT1 = 16'hf555;
    defparam sub_2065_add_2_29.INJECT1_0 = "NO";
    defparam sub_2065_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27179), .COUT(n27180));
    defparam sub_2065_add_2_27.INIT0 = 16'hf555;
    defparam sub_2065_add_2_27.INIT1 = 16'hf555;
    defparam sub_2065_add_2_27.INJECT1_0 = "NO";
    defparam sub_2065_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27178), .COUT(n27179));
    defparam sub_2065_add_2_25.INIT0 = 16'hf555;
    defparam sub_2065_add_2_25.INIT1 = 16'hf555;
    defparam sub_2065_add_2_25.INJECT1_0 = "NO";
    defparam sub_2065_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27177), .COUT(n27178));
    defparam sub_2065_add_2_23.INIT0 = 16'hf555;
    defparam sub_2065_add_2_23.INIT1 = 16'hf555;
    defparam sub_2065_add_2_23.INJECT1_0 = "NO";
    defparam sub_2065_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27176), .COUT(n27177));
    defparam sub_2065_add_2_21.INIT0 = 16'hf555;
    defparam sub_2065_add_2_21.INIT1 = 16'hf555;
    defparam sub_2065_add_2_21.INJECT1_0 = "NO";
    defparam sub_2065_add_2_21.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27579), .COUT(n27580), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2664_add_4_27.INJECT1_0 = "NO";
    defparam count_2664_add_4_27.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27175), .COUT(n27176));
    defparam sub_2065_add_2_19.INIT0 = 16'hf555;
    defparam sub_2065_add_2_19.INIT1 = 16'hf555;
    defparam sub_2065_add_2_19.INJECT1_0 = "NO";
    defparam sub_2065_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27174), .COUT(n27175));
    defparam sub_2065_add_2_17.INIT0 = 16'hf555;
    defparam sub_2065_add_2_17.INIT1 = 16'hf555;
    defparam sub_2065_add_2_17.INJECT1_0 = "NO";
    defparam sub_2065_add_2_17.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27578), .COUT(n27579), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2664_add_4_25.INJECT1_0 = "NO";
    defparam count_2664_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27577), .COUT(n27578), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2664_add_4_23.INJECT1_0 = "NO";
    defparam count_2664_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27576), .COUT(n27577), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2664_add_4_21.INJECT1_0 = "NO";
    defparam count_2664_add_4_21.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27173), .COUT(n27174));
    defparam sub_2065_add_2_15.INIT0 = 16'hf555;
    defparam sub_2065_add_2_15.INIT1 = 16'hf555;
    defparam sub_2065_add_2_15.INJECT1_0 = "NO";
    defparam sub_2065_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27172), .COUT(n27173));
    defparam sub_2065_add_2_13.INIT0 = 16'hf555;
    defparam sub_2065_add_2_13.INIT1 = 16'hf555;
    defparam sub_2065_add_2_13.INJECT1_0 = "NO";
    defparam sub_2065_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27171), .COUT(n27172));
    defparam sub_2065_add_2_11.INIT0 = 16'hf555;
    defparam sub_2065_add_2_11.INIT1 = 16'hf555;
    defparam sub_2065_add_2_11.INJECT1_0 = "NO";
    defparam sub_2065_add_2_11.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27575), .COUT(n27576), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2664_add_4_19.INJECT1_0 = "NO";
    defparam count_2664_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27574), .COUT(n27575), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2664_add_4_17.INJECT1_0 = "NO";
    defparam count_2664_add_4_17.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27170), .COUT(n27171));
    defparam sub_2065_add_2_9.INIT0 = 16'hf555;
    defparam sub_2065_add_2_9.INIT1 = 16'hf555;
    defparam sub_2065_add_2_9.INJECT1_0 = "NO";
    defparam sub_2065_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27169), .COUT(n27170));
    defparam sub_2065_add_2_7.INIT0 = 16'hf555;
    defparam sub_2065_add_2_7.INIT1 = 16'hf555;
    defparam sub_2065_add_2_7.INJECT1_0 = "NO";
    defparam sub_2065_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27168), .COUT(n27169));
    defparam sub_2065_add_2_5.INIT0 = 16'hf555;
    defparam sub_2065_add_2_5.INIT1 = 16'hf555;
    defparam sub_2065_add_2_5.INJECT1_0 = "NO";
    defparam sub_2065_add_2_5.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27573), .COUT(n27574), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2664_add_4_15.INJECT1_0 = "NO";
    defparam count_2664_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27572), .COUT(n27573), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2664_add_4_13.INJECT1_0 = "NO";
    defparam count_2664_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27571), .COUT(n27572), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2664_add_4_11.INJECT1_0 = "NO";
    defparam count_2664_add_4_11.INJECT1_1 = "NO";
    CCU2D sub_2065_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27167), .COUT(n27168));
    defparam sub_2065_add_2_3.INIT0 = 16'hf555;
    defparam sub_2065_add_2_3.INIT1 = 16'hf555;
    defparam sub_2065_add_2_3.INJECT1_0 = "NO";
    defparam sub_2065_add_2_3.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27570), .COUT(n27571), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2664_add_4_9.INJECT1_0 = "NO";
    defparam count_2664_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27569), .COUT(n27570), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2664_add_4_7.INJECT1_0 = "NO";
    defparam count_2664_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27568), .COUT(n27569), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2664_add_4_5.INJECT1_0 = "NO";
    defparam count_2664_add_4_5.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n32132), .CD(n16806), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D count_2664_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27567), .COUT(n27568), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2664_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2664_add_4_3.INJECT1_0 = "NO";
    defparam count_2664_add_4_3.INJECT1_1 = "NO";
    FD1S3IX count_2664__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i1.GSR = "ENABLED";
    CCU2D sub_2065_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27167));
    defparam sub_2065_add_2_1.INIT0 = 16'h0000;
    defparam sub_2065_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2065_add_2_1.INJECT1_0 = "NO";
    defparam sub_2065_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2664_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27567), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664_add_4_1.INIT0 = 16'hF000;
    defparam count_2664_add_4_1.INIT1 = 16'h0555;
    defparam count_2664_add_4_1.INJECT1_0 = "NO";
    defparam count_2664_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2664__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i2.GSR = "ENABLED";
    FD1S3IX count_2664__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i3.GSR = "ENABLED";
    FD1S3IX count_2664__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i4.GSR = "ENABLED";
    FD1S3IX count_2664__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i5.GSR = "ENABLED";
    FD1S3IX count_2664__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i6.GSR = "ENABLED";
    FD1S3IX count_2664__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i7.GSR = "ENABLED";
    FD1S3IX count_2664__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i8.GSR = "ENABLED";
    FD1S3IX count_2664__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i9.GSR = "ENABLED";
    FD1S3IX count_2664__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i10.GSR = "ENABLED";
    FD1S3IX count_2664__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i11.GSR = "ENABLED";
    FD1S3IX count_2664__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i12.GSR = "ENABLED";
    FD1S3IX count_2664__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i13.GSR = "ENABLED";
    FD1S3IX count_2664__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i14.GSR = "ENABLED";
    FD1S3IX count_2664__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i15.GSR = "ENABLED";
    FD1S3IX count_2664__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i16.GSR = "ENABLED";
    FD1S3IX count_2664__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i17.GSR = "ENABLED";
    FD1S3IX count_2664__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i18.GSR = "ENABLED";
    FD1S3IX count_2664__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i19.GSR = "ENABLED";
    FD1S3IX count_2664__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i20.GSR = "ENABLED";
    FD1S3IX count_2664__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i21.GSR = "ENABLED";
    FD1S3IX count_2664__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i22.GSR = "ENABLED";
    FD1S3IX count_2664__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i23.GSR = "ENABLED";
    FD1S3IX count_2664__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i24.GSR = "ENABLED";
    FD1S3IX count_2664__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i25.GSR = "ENABLED";
    FD1S3IX count_2664__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i26.GSR = "ENABLED";
    FD1S3IX count_2664__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i27.GSR = "ENABLED";
    FD1S3IX count_2664__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i28.GSR = "ENABLED";
    FD1S3IX count_2664__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i29.GSR = "ENABLED";
    FD1S3IX count_2664__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i30.GSR = "ENABLED";
    FD1S3IX count_2664__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n32132), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2664__i31.GSR = "ENABLED";
    LUT4 i1028_2_lut_rep_311 (.A(n8204), .B(n34065), .Z(n32132)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i1028_2_lut_rep_311.init = 16'heeee;
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27526), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27525), .COUT(n27526), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27524), .COUT(n27525), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    LUT4 i10114_2_lut_3_lut (.A(n8204), .B(n34065), .C(n8238), .Z(n16806)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i10114_2_lut_3_lut.init = 16'he0e0;
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27523), .COUT(n27524), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27522), .COUT(n27523), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27521), .COUT(n27522), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27520), .COUT(n27521), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27519), .COUT(n27520), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27518), .COUT(n27519), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27517), .COUT(n27518), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27516), .COUT(n27517), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27515), .COUT(n27516), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27514), .COUT(n27515), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27513), .COUT(n27514), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27512), .COUT(n27513), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module ClockDivider_U10
//

module ClockDivider_U10 (n34065, n7822, n30615, n28233, n30621, n28222, 
            n30619, n28231, debug_c_c, n241, n30482, n13605, GND_net, 
            n32135, n30472, n13974, n30613, n28234, n30623, n28140, 
            n30617, n28232, n30470, n13975, n30465, n13976, n30463, 
            n13977, n30474, n32134) /* synthesis syn_module_defined=1 */ ;
    input n34065;
    output n7822;
    input n30615;
    output n28233;
    input n30621;
    output n28222;
    input n30619;
    output n28231;
    input debug_c_c;
    input n241;
    input n30482;
    output n13605;
    input GND_net;
    output n32135;
    input n30472;
    output n13974;
    input n30613;
    output n28234;
    input n30623;
    output n28140;
    input n30617;
    output n28232;
    input n30470;
    output n13975;
    input n30465;
    output n13976;
    input n30463;
    output n13977;
    input n30474;
    output n32134;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire clk_255kHz;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    
    wire n2764;
    wire [31:0]n134;
    
    wire n7857, n27752, n27751, n27750, n27749, n27748, n27747, 
        n27746, n27745, n27744, n27743, n27742, n27741, n27740, 
        n27739, n27738, n27326, n27325, n27324, n27323, n27322, 
        n27321, n27320, n27319, n27414, n27413, n27412, n27411, 
        n27410, n27318, n27317, n27409, n27408, n27316, n27315, 
        n27407, n27406, n27314, n27405, n27404, n27313, n27312, 
        n27311, n27403, n27402, n27401, n27400, n27399;
    
    LUT4 i23214_2_lut_4_lut (.A(n34065), .B(clk_255kHz), .C(n7822), .D(n30615), 
         .Z(n28233)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23214_2_lut_4_lut.init = 16'h1000;
    LUT4 i23220_2_lut_4_lut (.A(n34065), .B(clk_255kHz), .C(n7822), .D(n30621), 
         .Z(n28222)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23220_2_lut_4_lut.init = 16'h1000;
    LUT4 i23218_2_lut_4_lut (.A(n34065), .B(clk_255kHz), .C(n7822), .D(n30619), 
         .Z(n28231)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23218_2_lut_4_lut.init = 16'h1000;
    FD1S3AX clk_o_22 (.D(n241), .CK(debug_c_c), .Q(clk_255kHz)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=540, LSE_RLINE=543 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    FD1S3IX count_2659__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2764), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i0.GSR = "ENABLED";
    LUT4 i962_2_lut (.A(n7857), .B(n34065), .Z(n2764)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i962_2_lut.init = 16'heeee;
    LUT4 i23081_2_lut_4_lut (.A(n34065), .B(clk_255kHz), .C(n7822), .D(n30482), 
         .Z(n13605)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23081_2_lut_4_lut.init = 16'h1000;
    CCU2D add_20293_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27752), 
          .S1(n7822));
    defparam add_20293_32.INIT0 = 16'h5555;
    defparam add_20293_32.INIT1 = 16'h0000;
    defparam add_20293_32.INJECT1_0 = "NO";
    defparam add_20293_32.INJECT1_1 = "NO";
    CCU2D add_20293_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27751), .COUT(n27752));
    defparam add_20293_30.INIT0 = 16'h5555;
    defparam add_20293_30.INIT1 = 16'h5555;
    defparam add_20293_30.INJECT1_0 = "NO";
    defparam add_20293_30.INJECT1_1 = "NO";
    CCU2D add_20293_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27750), .COUT(n27751));
    defparam add_20293_28.INIT0 = 16'h5555;
    defparam add_20293_28.INIT1 = 16'h5555;
    defparam add_20293_28.INJECT1_0 = "NO";
    defparam add_20293_28.INJECT1_1 = "NO";
    CCU2D add_20293_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27749), .COUT(n27750));
    defparam add_20293_26.INIT0 = 16'h5555;
    defparam add_20293_26.INIT1 = 16'h5555;
    defparam add_20293_26.INJECT1_0 = "NO";
    defparam add_20293_26.INJECT1_1 = "NO";
    CCU2D add_20293_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27748), .COUT(n27749));
    defparam add_20293_24.INIT0 = 16'h5555;
    defparam add_20293_24.INIT1 = 16'h5555;
    defparam add_20293_24.INJECT1_0 = "NO";
    defparam add_20293_24.INJECT1_1 = "NO";
    CCU2D add_20293_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27747), .COUT(n27748));
    defparam add_20293_22.INIT0 = 16'h5555;
    defparam add_20293_22.INIT1 = 16'h5555;
    defparam add_20293_22.INJECT1_0 = "NO";
    defparam add_20293_22.INJECT1_1 = "NO";
    CCU2D add_20293_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27746), .COUT(n27747));
    defparam add_20293_20.INIT0 = 16'h5555;
    defparam add_20293_20.INIT1 = 16'h5555;
    defparam add_20293_20.INJECT1_0 = "NO";
    defparam add_20293_20.INJECT1_1 = "NO";
    CCU2D add_20293_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27745), .COUT(n27746));
    defparam add_20293_18.INIT0 = 16'h5555;
    defparam add_20293_18.INIT1 = 16'h5555;
    defparam add_20293_18.INJECT1_0 = "NO";
    defparam add_20293_18.INJECT1_1 = "NO";
    CCU2D add_20293_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27744), .COUT(n27745));
    defparam add_20293_16.INIT0 = 16'h5555;
    defparam add_20293_16.INIT1 = 16'h5555;
    defparam add_20293_16.INJECT1_0 = "NO";
    defparam add_20293_16.INJECT1_1 = "NO";
    CCU2D add_20293_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27743), .COUT(n27744));
    defparam add_20293_14.INIT0 = 16'h5555;
    defparam add_20293_14.INIT1 = 16'h5555;
    defparam add_20293_14.INJECT1_0 = "NO";
    defparam add_20293_14.INJECT1_1 = "NO";
    CCU2D add_20293_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27742), .COUT(n27743));
    defparam add_20293_12.INIT0 = 16'h5555;
    defparam add_20293_12.INIT1 = 16'h5555;
    defparam add_20293_12.INJECT1_0 = "NO";
    defparam add_20293_12.INJECT1_1 = "NO";
    CCU2D add_20293_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27741), .COUT(n27742));
    defparam add_20293_10.INIT0 = 16'h5555;
    defparam add_20293_10.INIT1 = 16'h5555;
    defparam add_20293_10.INJECT1_0 = "NO";
    defparam add_20293_10.INJECT1_1 = "NO";
    CCU2D add_20293_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27740), 
          .COUT(n27741));
    defparam add_20293_8.INIT0 = 16'h5555;
    defparam add_20293_8.INIT1 = 16'h5555;
    defparam add_20293_8.INJECT1_0 = "NO";
    defparam add_20293_8.INJECT1_1 = "NO";
    CCU2D add_20293_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27739), 
          .COUT(n27740));
    defparam add_20293_6.INIT0 = 16'h5555;
    defparam add_20293_6.INIT1 = 16'h5555;
    defparam add_20293_6.INJECT1_0 = "NO";
    defparam add_20293_6.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_314 (.A(n34065), .B(clk_255kHz), .C(n7822), .Z(n32135)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i2_3_lut_rep_314.init = 16'h1010;
    CCU2D add_20293_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27738), 
          .COUT(n27739));
    defparam add_20293_4.INIT0 = 16'h5555;
    defparam add_20293_4.INIT1 = 16'h5aaa;
    defparam add_20293_4.INJECT1_0 = "NO";
    defparam add_20293_4.INJECT1_1 = "NO";
    CCU2D add_20293_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27738));
    defparam add_20293_2.INIT0 = 16'h7000;
    defparam add_20293_2.INIT1 = 16'h5aaa;
    defparam add_20293_2.INJECT1_0 = "NO";
    defparam add_20293_2.INJECT1_1 = "NO";
    FD1S3IX count_2659__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2764), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i1.GSR = "ENABLED";
    FD1S3IX count_2659__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2764), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i2.GSR = "ENABLED";
    FD1S3IX count_2659__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2764), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i3.GSR = "ENABLED";
    FD1S3IX count_2659__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2764), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i4.GSR = "ENABLED";
    FD1S3IX count_2659__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2764), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i5.GSR = "ENABLED";
    FD1S3IX count_2659__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2764), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i6.GSR = "ENABLED";
    FD1S3IX count_2659__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2764), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i7.GSR = "ENABLED";
    FD1S3IX count_2659__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2764), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i8.GSR = "ENABLED";
    FD1S3IX count_2659__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2764), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i9.GSR = "ENABLED";
    FD1S3IX count_2659__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i10.GSR = "ENABLED";
    FD1S3IX count_2659__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i11.GSR = "ENABLED";
    FD1S3IX count_2659__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i12.GSR = "ENABLED";
    FD1S3IX count_2659__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i13.GSR = "ENABLED";
    FD1S3IX count_2659__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i14.GSR = "ENABLED";
    FD1S3IX count_2659__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i15.GSR = "ENABLED";
    FD1S3IX count_2659__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i16.GSR = "ENABLED";
    FD1S3IX count_2659__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i17.GSR = "ENABLED";
    FD1S3IX count_2659__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i18.GSR = "ENABLED";
    FD1S3IX count_2659__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i19.GSR = "ENABLED";
    FD1S3IX count_2659__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i20.GSR = "ENABLED";
    FD1S3IX count_2659__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i21.GSR = "ENABLED";
    FD1S3IX count_2659__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i22.GSR = "ENABLED";
    FD1S3IX count_2659__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i23.GSR = "ENABLED";
    FD1S3IX count_2659__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i24.GSR = "ENABLED";
    FD1S3IX count_2659__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i25.GSR = "ENABLED";
    FD1S3IX count_2659__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i26.GSR = "ENABLED";
    FD1S3IX count_2659__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i27.GSR = "ENABLED";
    FD1S3IX count_2659__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i28.GSR = "ENABLED";
    FD1S3IX count_2659__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i29.GSR = "ENABLED";
    FD1S3IX count_2659__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i30.GSR = "ENABLED";
    FD1S3IX count_2659__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2764), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659__i31.GSR = "ENABLED";
    LUT4 i23071_2_lut_4_lut (.A(n34065), .B(clk_255kHz), .C(n7822), .D(n30472), 
         .Z(n13974)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23071_2_lut_4_lut.init = 16'h1000;
    LUT4 i23212_2_lut_4_lut (.A(n34065), .B(clk_255kHz), .C(n7822), .D(n30613), 
         .Z(n28234)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23212_2_lut_4_lut.init = 16'h1000;
    CCU2D sub_2047_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27326), .S0(n7857));
    defparam sub_2047_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2047_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2047_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2047_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27325), .COUT(n27326));
    defparam sub_2047_add_2_32.INIT0 = 16'h5555;
    defparam sub_2047_add_2_32.INIT1 = 16'h5555;
    defparam sub_2047_add_2_32.INJECT1_0 = "NO";
    defparam sub_2047_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27324), .COUT(n27325));
    defparam sub_2047_add_2_30.INIT0 = 16'h5555;
    defparam sub_2047_add_2_30.INIT1 = 16'h5555;
    defparam sub_2047_add_2_30.INJECT1_0 = "NO";
    defparam sub_2047_add_2_30.INJECT1_1 = "NO";
    LUT4 i23222_2_lut_4_lut (.A(n34065), .B(clk_255kHz), .C(n7822), .D(n30623), 
         .Z(n28140)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23222_2_lut_4_lut.init = 16'h1000;
    CCU2D sub_2047_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27323), .COUT(n27324));
    defparam sub_2047_add_2_28.INIT0 = 16'h5555;
    defparam sub_2047_add_2_28.INIT1 = 16'h5555;
    defparam sub_2047_add_2_28.INJECT1_0 = "NO";
    defparam sub_2047_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27322), .COUT(n27323));
    defparam sub_2047_add_2_26.INIT0 = 16'h5555;
    defparam sub_2047_add_2_26.INIT1 = 16'h5555;
    defparam sub_2047_add_2_26.INJECT1_0 = "NO";
    defparam sub_2047_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27321), .COUT(n27322));
    defparam sub_2047_add_2_24.INIT0 = 16'h5555;
    defparam sub_2047_add_2_24.INIT1 = 16'h5555;
    defparam sub_2047_add_2_24.INJECT1_0 = "NO";
    defparam sub_2047_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27320), .COUT(n27321));
    defparam sub_2047_add_2_22.INIT0 = 16'h5555;
    defparam sub_2047_add_2_22.INIT1 = 16'h5555;
    defparam sub_2047_add_2_22.INJECT1_0 = "NO";
    defparam sub_2047_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27319), .COUT(n27320));
    defparam sub_2047_add_2_20.INIT0 = 16'h5555;
    defparam sub_2047_add_2_20.INIT1 = 16'h5555;
    defparam sub_2047_add_2_20.INJECT1_0 = "NO";
    defparam sub_2047_add_2_20.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27414), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_33.INIT1 = 16'h0000;
    defparam count_2659_add_4_33.INJECT1_0 = "NO";
    defparam count_2659_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27413), .COUT(n27414), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2659_add_4_31.INJECT1_0 = "NO";
    defparam count_2659_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27412), .COUT(n27413), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2659_add_4_29.INJECT1_0 = "NO";
    defparam count_2659_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27411), .COUT(n27412), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2659_add_4_27.INJECT1_0 = "NO";
    defparam count_2659_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27410), .COUT(n27411), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2659_add_4_25.INJECT1_0 = "NO";
    defparam count_2659_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27318), .COUT(n27319));
    defparam sub_2047_add_2_18.INIT0 = 16'h5555;
    defparam sub_2047_add_2_18.INIT1 = 16'h5555;
    defparam sub_2047_add_2_18.INJECT1_0 = "NO";
    defparam sub_2047_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27317), .COUT(n27318));
    defparam sub_2047_add_2_16.INIT0 = 16'h5555;
    defparam sub_2047_add_2_16.INIT1 = 16'h5555;
    defparam sub_2047_add_2_16.INJECT1_0 = "NO";
    defparam sub_2047_add_2_16.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27409), .COUT(n27410), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2659_add_4_23.INJECT1_0 = "NO";
    defparam count_2659_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27408), .COUT(n27409), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2659_add_4_21.INJECT1_0 = "NO";
    defparam count_2659_add_4_21.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27316), .COUT(n27317));
    defparam sub_2047_add_2_14.INIT0 = 16'h5555;
    defparam sub_2047_add_2_14.INIT1 = 16'h5555;
    defparam sub_2047_add_2_14.INJECT1_0 = "NO";
    defparam sub_2047_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27315), .COUT(n27316));
    defparam sub_2047_add_2_12.INIT0 = 16'h5555;
    defparam sub_2047_add_2_12.INIT1 = 16'h5555;
    defparam sub_2047_add_2_12.INJECT1_0 = "NO";
    defparam sub_2047_add_2_12.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27407), .COUT(n27408), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2659_add_4_19.INJECT1_0 = "NO";
    defparam count_2659_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27406), .COUT(n27407), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2659_add_4_17.INJECT1_0 = "NO";
    defparam count_2659_add_4_17.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27314), .COUT(n27315));
    defparam sub_2047_add_2_10.INIT0 = 16'h5555;
    defparam sub_2047_add_2_10.INIT1 = 16'h5555;
    defparam sub_2047_add_2_10.INJECT1_0 = "NO";
    defparam sub_2047_add_2_10.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27405), .COUT(n27406), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2659_add_4_15.INJECT1_0 = "NO";
    defparam count_2659_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27404), .COUT(n27405), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2659_add_4_13.INJECT1_0 = "NO";
    defparam count_2659_add_4_13.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27313), .COUT(n27314));
    defparam sub_2047_add_2_8.INIT0 = 16'h5555;
    defparam sub_2047_add_2_8.INIT1 = 16'h5555;
    defparam sub_2047_add_2_8.INJECT1_0 = "NO";
    defparam sub_2047_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27312), .COUT(n27313));
    defparam sub_2047_add_2_6.INIT0 = 16'h5555;
    defparam sub_2047_add_2_6.INIT1 = 16'h5aaa;
    defparam sub_2047_add_2_6.INJECT1_0 = "NO";
    defparam sub_2047_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27311), .COUT(n27312));
    defparam sub_2047_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2047_add_2_4.INIT1 = 16'h5aaa;
    defparam sub_2047_add_2_4.INJECT1_0 = "NO";
    defparam sub_2047_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_2047_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27311));
    defparam sub_2047_add_2_2.INIT0 = 16'h0000;
    defparam sub_2047_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2047_add_2_2.INJECT1_0 = "NO";
    defparam sub_2047_add_2_2.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27403), .COUT(n27404), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2659_add_4_11.INJECT1_0 = "NO";
    defparam count_2659_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27402), .COUT(n27403), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2659_add_4_9.INJECT1_0 = "NO";
    defparam count_2659_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27401), .COUT(n27402), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2659_add_4_7.INJECT1_0 = "NO";
    defparam count_2659_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27400), .COUT(n27401), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2659_add_4_5.INJECT1_0 = "NO";
    defparam count_2659_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27399), .COUT(n27400), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2659_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2659_add_4_3.INJECT1_0 = "NO";
    defparam count_2659_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2659_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27399), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2659_add_4_1.INIT0 = 16'hF000;
    defparam count_2659_add_4_1.INIT1 = 16'h0555;
    defparam count_2659_add_4_1.INJECT1_0 = "NO";
    defparam count_2659_add_4_1.INJECT1_1 = "NO";
    LUT4 i23216_2_lut_4_lut (.A(n34065), .B(clk_255kHz), .C(n7822), .D(n30617), 
         .Z(n28232)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23216_2_lut_4_lut.init = 16'h1000;
    LUT4 i23069_2_lut_4_lut (.A(n34065), .B(clk_255kHz), .C(n7822), .D(n30470), 
         .Z(n13975)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23069_2_lut_4_lut.init = 16'h1000;
    LUT4 i23064_2_lut_4_lut (.A(n34065), .B(clk_255kHz), .C(n7822), .D(n30465), 
         .Z(n13976)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23064_2_lut_4_lut.init = 16'h1000;
    LUT4 i23062_2_lut_4_lut (.A(n34065), .B(clk_255kHz), .C(n7822), .D(n30463), 
         .Z(n13977)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23062_2_lut_4_lut.init = 16'h1000;
    LUT4 i23073_2_lut_rep_313_4_lut (.A(n34065), .B(clk_255kHz), .C(n7822), 
         .D(n30474), .Z(n32134)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i23073_2_lut_rep_313_4_lut.init = 16'h1000;
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b010000) 
//

module \ArmPeripheral(axis_haddr=8'b010000)  (debug_c_c, n34070, n34069, 
            \register_addr[0] , VCC_net, GND_net, Stepper_Y_nFault_c, 
            n34066, \read_size[0] , n2776, n29713, Stepper_Y_M0_c_0, 
            n13899, n579, prev_step_clk, step_clk, n13885, prev_select, 
            n32163, read_value, Stepper_Y_Step_c, n32140, n34067, 
            databus, n34071, n608, \control_reg[7] , n13576, Stepper_Y_En_c, 
            Stepper_Y_Dir_c, Stepper_Y_M2_c_2, Stepper_Y_M1_c_1, n4034, 
            \read_size[2] , n28426, n34068, \register_addr[1] , limit_c_1, 
            n34065, n32, n22, n32144, n8576, n28049) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n34070;
    input n34069;
    input \register_addr[0] ;
    input VCC_net;
    input GND_net;
    input Stepper_Y_nFault_c;
    input n34066;
    output \read_size[0] ;
    input n2776;
    input n29713;
    output Stepper_Y_M0_c_0;
    input n13899;
    input n579;
    output prev_step_clk;
    output step_clk;
    input n13885;
    output prev_select;
    input n32163;
    output [31:0]read_value;
    output Stepper_Y_Step_c;
    input n32140;
    input n34067;
    input [31:0]databus;
    input n34071;
    input n608;
    output \control_reg[7] ;
    input n13576;
    output Stepper_Y_En_c;
    output Stepper_Y_Dir_c;
    output Stepper_Y_M2_c_2;
    output Stepper_Y_M1_c_1;
    input n4034;
    output \read_size[2] ;
    input n28426;
    input n34068;
    input \register_addr[1] ;
    input limit_c_1;
    input n34065;
    input n32;
    input n22;
    input n32144;
    input n8576;
    output n28049;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n4035;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]n6683;
    
    wire fault_latched, limit_latched, n30348, n30349, n182, prev_limit_latched, 
        n30350;
    wire [31:0]n100;
    
    wire n30410, n30368, int_step;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n11186;
    wire [31:0]n224;
    
    wire n30408, n30409, n30366, n30367, n27446, n27445, n27444, 
        n27443, n27442, n27441, n27440, n27439, n27438, n27437, 
        n27436, n27435, n27434, n27433, n27432, n27431;
    wire [7:0]n8575;
    
    wire n49, n62_adj_557, n58_adj_558, n50_adj_559, n41, n60_adj_560, 
        n54_adj_561, n42_adj_562, n52_adj_563, n38_adj_564, n56_adj_565, 
        n46_adj_566;
    
    FD1S3IX steps_reg__i13 (.D(n4035[13]), .CK(debug_c_c), .CD(n34070), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n4035[12]), .CK(debug_c_c), .CD(n34070), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n4035[11]), .CK(debug_c_c), .CD(n34070), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n4035[10]), .CK(debug_c_c), .CD(n34070), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n4035[9]), .CK(debug_c_c), .CD(n34070), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n4035[8]), .CK(debug_c_c), .CD(n34070), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n4035[7]), .CK(debug_c_c), .CD(n34070), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n4035[6]), .CK(debug_c_c), .CD(n34070), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n4035[5]), .CK(debug_c_c), .CD(n34070), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n4035[4]), .CK(debug_c_c), .CD(n34069), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n4035[3]), .CK(debug_c_c), .CD(n34069), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n4035[2]), .CK(debug_c_c), .CD(n34069), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n4035[1]), .CK(debug_c_c), .CD(n34069), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 mux_1938_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n6683[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1938_i8_3_lut.init = 16'hcaca;
    IFS1P3DX fault_latched_178 (.D(Stepper_Y_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n4035[0]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n29713), .SP(n2776), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    LUT4 i22845_3_lut (.A(Stepper_Y_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n30348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22845_3_lut.init = 16'hcaca;
    LUT4 i22846_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n30349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22846_3_lut.init = 16'hcaca;
    FD1P3AX control_reg_i1 (.D(n579), .SP(n13899), .CK(debug_c_c), .Q(Stepper_Y_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n13885), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n32163), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n30350), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n100[26]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n100[23]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n100[20]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n100[7]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30410), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30368), .SP(n2776), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_Y_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n32140), .PD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n32140), .PD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n32140), .PD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n32140), .PD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n32140), .PD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n32140), .PD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n32140), .PD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n13885), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n13576), .CD(n11186), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n13576), .PD(n34067), 
            .CK(debug_c_c), .Q(Stepper_Y_En_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n13576), .PD(n34067), 
            .CK(debug_c_c), .Q(Stepper_Y_Dir_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n13899), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n13576), .PD(n34067), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n13576), .CD(n34067), 
            .CK(debug_c_c), .Q(Stepper_Y_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n13576), .PD(n34067), 
            .CK(debug_c_c), .Q(Stepper_Y_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    LUT4 mux_1587_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n4034), 
         .Z(n4035[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i14_3_lut.init = 16'hcaca;
    FD1P3AX read_size__i2 (.D(n28426), .SP(n2776), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n4035[31]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n4035[30]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n4035[29]), .CK(debug_c_c), .CD(n34071), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n4035[28]), .CK(debug_c_c), .CD(n34071), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n4035[27]), .CK(debug_c_c), .CD(n34071), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n4035[26]), .CK(debug_c_c), .CD(n34071), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n4035[25]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n4035[24]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n4035[23]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n4035[22]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n4035[21]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n4035[20]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n4035[19]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n4035[18]), .CK(debug_c_c), .CD(n34071), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n4035[17]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n4035[16]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n4035[15]), .CK(debug_c_c), .CD(n34071), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    PFUMX i22907 (.BLUT(n30408), .ALUT(n30409), .C0(\register_addr[0] ), 
          .Z(n30410));
    LUT4 mux_1587_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n4034), 
         .Z(n4035[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n4034), 
         .Z(n4035[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n4034), 
         .Z(n4035[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n4034), .Z(n4035[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n4034), .Z(n4035[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n4034), .Z(n4035[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n4034), .Z(n4035[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n4034), .Z(n4035[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n4034), .Z(n4035[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i10_3_lut.init = 16'hcaca;
    LUT4 i15272_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15272_4_lut.init = 16'hc088;
    LUT4 i15273_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15273_4_lut.init = 16'hc088;
    LUT4 i15274_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15274_4_lut.init = 16'hc088;
    LUT4 i15275_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15275_4_lut.init = 16'hc088;
    LUT4 i15276_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15276_4_lut.init = 16'hc088;
    LUT4 i15277_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n100[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15277_4_lut.init = 16'hc088;
    LUT4 i15278_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15278_4_lut.init = 16'hc088;
    LUT4 i15279_4_lut (.A(div_factor_reg[24]), .B(\register_addr[1] ), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15279_4_lut.init = 16'hc088;
    LUT4 i15280_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n100[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15280_4_lut.init = 16'hc088;
    LUT4 i15281_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15281_4_lut.init = 16'hc088;
    LUT4 i15282_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15282_4_lut.init = 16'hc088;
    LUT4 i15283_4_lut (.A(div_factor_reg[20]), .B(\register_addr[1] ), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n100[20])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15283_4_lut.init = 16'hc088;
    LUT4 i15284_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15284_4_lut.init = 16'hc088;
    LUT4 i15285_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15285_4_lut.init = 16'hc088;
    LUT4 i15286_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15286_4_lut.init = 16'hc088;
    LUT4 i15287_4_lut (.A(div_factor_reg[16]), .B(\register_addr[1] ), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n100[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15287_4_lut.init = 16'hc088;
    LUT4 i15288_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15288_4_lut.init = 16'hc088;
    LUT4 i15289_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15289_4_lut.init = 16'hc088;
    LUT4 i15290_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15290_4_lut.init = 16'hc088;
    LUT4 i15291_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15291_4_lut.init = 16'hc088;
    LUT4 i15292_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15292_4_lut.init = 16'hc088;
    LUT4 i15293_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15293_4_lut.init = 16'hc088;
    LUT4 i118_1_lut (.A(limit_c_1), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i15294_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15294_4_lut.init = 16'hc088;
    LUT4 i15295_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15295_4_lut.init = 16'hc088;
    LUT4 mux_1587_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n4034), .Z(n4035[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n4034), 
         .Z(n4035[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i12_3_lut.init = 16'hcaca;
    PFUMX i22847 (.BLUT(n30348), .ALUT(n30349), .C0(\register_addr[1] ), 
          .Z(n30350));
    LUT4 mux_1587_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n4034), .Z(n4035[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i7_3_lut.init = 16'hcaca;
    LUT4 i4470_3_lut (.A(prev_limit_latched), .B(n34065), .C(limit_latched), 
         .Z(n11186)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i4470_3_lut.init = 16'hdcdc;
    LUT4 i22863_3_lut (.A(Stepper_Y_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n30366)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22863_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i14 (.D(n4035[14]), .CK(debug_c_c), .CD(n34070), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    LUT4 i22864_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n30367)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22864_3_lut.init = 16'hcaca;
    PFUMX i22865 (.BLUT(n30366), .ALUT(n30367), .C0(\register_addr[1] ), 
          .Z(n30368));
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27446), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27445), .COUT(n27446), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27444), .COUT(n27445), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27443), .COUT(n27444), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27442), .COUT(n27443), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27441), .COUT(n27442), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27440), .COUT(n27441), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27439), .COUT(n27440), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27438), .COUT(n27439), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27437), .COUT(n27438), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n13885), .CD(n34067), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n13885), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n13885), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n13885), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n13885), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n13885), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n13885), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n13885), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n13885), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n13885), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n13885), .CD(n34070), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n13885), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n13885), .CD(n34070), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n13885), .CD(n34070), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n13885), .CD(n34070), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27436), .COUT(n27437), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n13885), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n13885), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n13885), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n13885), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n13885), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n13885), .CD(n34070), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n13885), .CD(n34070), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n13885), .CD(n34070), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=595, LSE_RLINE=608 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27435), .COUT(n27436), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27434), .COUT(n27435), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27433), .COUT(n27434), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27432), .COUT(n27433), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27431), .COUT(n27432), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n27431), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    FD1P3AX int_step_182 (.D(n32144), .SP(n22), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 mux_1587_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n4034), .Z(n4035[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n4034), 
         .Z(n4035[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n4034), 
         .Z(n4035[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n4034), 
         .Z(n4035[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n4034), 
         .Z(n4035[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n4034), 
         .Z(n4035[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n4034), 
         .Z(n4035[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n4034), 
         .Z(n4035[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n4034), 
         .Z(n4035[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n4034), 
         .Z(n4035[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n4034), 
         .Z(n4035[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n4034), 
         .Z(n4035[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n4034), 
         .Z(n4035[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n4034), 
         .Z(n4035[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n4034), 
         .Z(n4035[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n4034), 
         .Z(n4035[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n4034), 
         .Z(n4035[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1587_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n4034), 
         .Z(n4035[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i16_3_lut.init = 16'hcaca;
    PFUMX mux_1942_i4 (.BLUT(n8575[3]), .ALUT(n6683[3]), .C0(\register_addr[1] ), 
          .Z(n100[3]));
    PFUMX mux_1942_i5 (.BLUT(n8575[4]), .ALUT(n6683[4]), .C0(\register_addr[1] ), 
          .Z(n100[4]));
    PFUMX mux_1942_i6 (.BLUT(n8575[5]), .ALUT(n6683[5]), .C0(\register_addr[1] ), 
          .Z(n100[5]));
    PFUMX mux_1942_i7 (.BLUT(n8575[6]), .ALUT(n6683[6]), .C0(\register_addr[1] ), 
          .Z(n100[6]));
    PFUMX mux_1942_i8 (.BLUT(n8576), .ALUT(n6683[7]), .C0(\register_addr[1] ), 
          .Z(n100[7]));
    LUT4 i22905_3_lut (.A(Stepper_Y_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n30408)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22905_3_lut.init = 16'hcaca;
    LUT4 i22906_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n30409)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22906_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62_adj_557), .C(n58_adj_558), .D(n50_adj_559), 
         .Z(n28049)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[0]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60_adj_560), .C(n54_adj_561), .D(n42_adj_562), 
         .Z(n62_adj_557)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52_adj_563), .C(n38_adj_564), 
         .D(steps_reg[18]), .Z(n58_adj_558)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50_adj_559)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[7]), .B(steps_reg[9]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[26]), .B(n56_adj_565), .C(n46_adj_566), 
         .D(steps_reg[29]), .Z(n60_adj_560)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 mux_1587_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n4034), .Z(n4035[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1587_i6_3_lut.init = 16'hcaca;
    LUT4 i22_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[25]), .Z(n54_adj_561)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n42_adj_562)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[10]), .B(steps_reg[22]), .C(steps_reg[20]), 
         .D(steps_reg[3]), .Z(n56_adj_565)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[5]), .B(steps_reg[6]), .Z(n46_adj_566)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[28]), .C(steps_reg[13]), 
         .D(steps_reg[30]), .Z(n52_adj_563)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[2]), .B(steps_reg[8]), .Z(n38_adj_564)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i15319_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n8575[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15319_2_lut.init = 16'h2222;
    LUT4 mux_1938_i4_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), .C(\register_addr[0] ), 
         .Z(n6683[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1938_i4_3_lut.init = 16'hcaca;
    LUT4 i15318_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n8575[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15318_2_lut.init = 16'h2222;
    LUT4 mux_1938_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n6683[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1938_i5_3_lut.init = 16'hcaca;
    LUT4 i15317_2_lut (.A(Stepper_Y_Dir_c), .B(\register_addr[0] ), .Z(n8575[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15317_2_lut.init = 16'h2222;
    LUT4 mux_1938_i6_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), .C(\register_addr[0] ), 
         .Z(n6683[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1938_i6_3_lut.init = 16'hcaca;
    LUT4 i15316_2_lut (.A(Stepper_Y_En_c), .B(\register_addr[0] ), .Z(n8575[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15316_2_lut.init = 16'h2222;
    LUT4 mux_1938_i7_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n6683[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1938_i7_3_lut.init = 16'hcaca;
    ClockDivider_U7 step_clk_gen (.div_factor_reg({div_factor_reg}), .GND_net(GND_net), 
            .step_clk(step_clk), .debug_c_c(debug_c_c), .n34071(n34071), 
            .n34065(n34065)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U7
//

module ClockDivider_U7 (div_factor_reg, GND_net, step_clk, debug_c_c, 
            n34071, n34065) /* synthesis syn_module_defined=1 */ ;
    input [31:0]div_factor_reg;
    input GND_net;
    output step_clk;
    input debug_c_c;
    input n34071;
    input n34065;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27222, n27223, n27221, n27220, n27219, n27510;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    wire [31:0]n40;
    
    wire n27509, n27218, n27508, n27507, n27217, n27506, n27505, 
        n27504, n27216, n27503, n27502, n27501, n27500, n27499, 
        n27498, n27497, n27215, n27496, n27495, n8065;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    
    wire n32130;
    wire [31:0]n134;
    
    wire n16775, n27262, n27261, n27260, n27259, n27258, n27257, 
        n27256, n27255, n27254, n27253, n27252, n27251, n27250, 
        n27249, n27248, n27247, n27246, n8100, n27245, n27244, 
        n27243, n27242, n27241, n27240, n27239, n27238, n27237, 
        n27236, n27235, n27234, n27694, n27693, n27233, n27692, 
        n27691, n27690, n27232, n27231, n27689, n27688, n27687, 
        n27686, n27685, n27684, n27683, n27682, n27681, n27680, 
        n27679, n27230, n8134, n27229, n27228, n27227, n27226, 
        n27225, n27224;
    
    CCU2D sub_2060_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27222), .COUT(n27223));
    defparam sub_2060_add_2_17.INIT0 = 16'hf555;
    defparam sub_2060_add_2_17.INIT1 = 16'hf555;
    defparam sub_2060_add_2_17.INJECT1_0 = "NO";
    defparam sub_2060_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2060_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27221), .COUT(n27222));
    defparam sub_2060_add_2_15.INIT0 = 16'hf555;
    defparam sub_2060_add_2_15.INIT1 = 16'hf555;
    defparam sub_2060_add_2_15.INJECT1_0 = "NO";
    defparam sub_2060_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2060_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27220), .COUT(n27221));
    defparam sub_2060_add_2_13.INIT0 = 16'hf555;
    defparam sub_2060_add_2_13.INIT1 = 16'hf555;
    defparam sub_2060_add_2_13.INJECT1_0 = "NO";
    defparam sub_2060_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2060_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27219), .COUT(n27220));
    defparam sub_2060_add_2_11.INIT0 = 16'hf555;
    defparam sub_2060_add_2_11.INIT1 = 16'hf555;
    defparam sub_2060_add_2_11.INJECT1_0 = "NO";
    defparam sub_2060_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27510), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27509), .COUT(n27510), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2060_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27218), .COUT(n27219));
    defparam sub_2060_add_2_9.INIT0 = 16'hf555;
    defparam sub_2060_add_2_9.INIT1 = 16'hf555;
    defparam sub_2060_add_2_9.INJECT1_0 = "NO";
    defparam sub_2060_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27508), .COUT(n27509), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27507), .COUT(n27508), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2060_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27217), .COUT(n27218));
    defparam sub_2060_add_2_7.INIT0 = 16'hf555;
    defparam sub_2060_add_2_7.INIT1 = 16'hf555;
    defparam sub_2060_add_2_7.INJECT1_0 = "NO";
    defparam sub_2060_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27506), .COUT(n27507), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27505), .COUT(n27506), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27504), .COUT(n27505), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2060_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27216), .COUT(n27217));
    defparam sub_2060_add_2_5.INIT0 = 16'hf555;
    defparam sub_2060_add_2_5.INIT1 = 16'hf555;
    defparam sub_2060_add_2_5.INJECT1_0 = "NO";
    defparam sub_2060_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27503), .COUT(n27504), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27502), .COUT(n27503), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27501), .COUT(n27502), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27500), .COUT(n27501), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27499), .COUT(n27500), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27498), .COUT(n27499), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27497), .COUT(n27498), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2060_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27215), .COUT(n27216));
    defparam sub_2060_add_2_3.INIT0 = 16'hf555;
    defparam sub_2060_add_2_3.INIT1 = 16'hf555;
    defparam sub_2060_add_2_3.INJECT1_0 = "NO";
    defparam sub_2060_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2060_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27215));
    defparam sub_2060_add_2_1.INIT0 = 16'h0000;
    defparam sub_2060_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2060_add_2_1.INJECT1_0 = "NO";
    defparam sub_2060_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27496), .COUT(n27497), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27495), .COUT(n27496), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27495), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n8065), .CK(debug_c_c), .CD(n34071), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    FD1S3IX count_2663__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i0.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n32130), .PD(n16775), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_2057_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27262), .S1(n8065));
    defparam sub_2057_add_2_33.INIT0 = 16'h5555;
    defparam sub_2057_add_2_33.INIT1 = 16'h0000;
    defparam sub_2057_add_2_33.INJECT1_0 = "NO";
    defparam sub_2057_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27261), .COUT(n27262));
    defparam sub_2057_add_2_31.INIT0 = 16'h5999;
    defparam sub_2057_add_2_31.INIT1 = 16'h5999;
    defparam sub_2057_add_2_31.INJECT1_0 = "NO";
    defparam sub_2057_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27260), .COUT(n27261));
    defparam sub_2057_add_2_29.INIT0 = 16'h5999;
    defparam sub_2057_add_2_29.INIT1 = 16'h5999;
    defparam sub_2057_add_2_29.INJECT1_0 = "NO";
    defparam sub_2057_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27259), .COUT(n27260));
    defparam sub_2057_add_2_27.INIT0 = 16'h5999;
    defparam sub_2057_add_2_27.INIT1 = 16'h5999;
    defparam sub_2057_add_2_27.INJECT1_0 = "NO";
    defparam sub_2057_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27258), .COUT(n27259));
    defparam sub_2057_add_2_25.INIT0 = 16'h5999;
    defparam sub_2057_add_2_25.INIT1 = 16'h5999;
    defparam sub_2057_add_2_25.INJECT1_0 = "NO";
    defparam sub_2057_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27257), .COUT(n27258));
    defparam sub_2057_add_2_23.INIT0 = 16'h5999;
    defparam sub_2057_add_2_23.INIT1 = 16'h5999;
    defparam sub_2057_add_2_23.INJECT1_0 = "NO";
    defparam sub_2057_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27256), .COUT(n27257));
    defparam sub_2057_add_2_21.INIT0 = 16'h5999;
    defparam sub_2057_add_2_21.INIT1 = 16'h5999;
    defparam sub_2057_add_2_21.INJECT1_0 = "NO";
    defparam sub_2057_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27255), .COUT(n27256));
    defparam sub_2057_add_2_19.INIT0 = 16'h5999;
    defparam sub_2057_add_2_19.INIT1 = 16'h5999;
    defparam sub_2057_add_2_19.INJECT1_0 = "NO";
    defparam sub_2057_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27254), .COUT(n27255));
    defparam sub_2057_add_2_17.INIT0 = 16'h5999;
    defparam sub_2057_add_2_17.INIT1 = 16'h5999;
    defparam sub_2057_add_2_17.INJECT1_0 = "NO";
    defparam sub_2057_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27253), .COUT(n27254));
    defparam sub_2057_add_2_15.INIT0 = 16'h5999;
    defparam sub_2057_add_2_15.INIT1 = 16'h5999;
    defparam sub_2057_add_2_15.INJECT1_0 = "NO";
    defparam sub_2057_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27252), .COUT(n27253));
    defparam sub_2057_add_2_13.INIT0 = 16'h5999;
    defparam sub_2057_add_2_13.INIT1 = 16'h5999;
    defparam sub_2057_add_2_13.INJECT1_0 = "NO";
    defparam sub_2057_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27251), .COUT(n27252));
    defparam sub_2057_add_2_11.INIT0 = 16'h5999;
    defparam sub_2057_add_2_11.INIT1 = 16'h5999;
    defparam sub_2057_add_2_11.INJECT1_0 = "NO";
    defparam sub_2057_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27250), .COUT(n27251));
    defparam sub_2057_add_2_9.INIT0 = 16'h5999;
    defparam sub_2057_add_2_9.INIT1 = 16'h5999;
    defparam sub_2057_add_2_9.INJECT1_0 = "NO";
    defparam sub_2057_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27249), .COUT(n27250));
    defparam sub_2057_add_2_7.INIT0 = 16'h5999;
    defparam sub_2057_add_2_7.INIT1 = 16'h5999;
    defparam sub_2057_add_2_7.INJECT1_0 = "NO";
    defparam sub_2057_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27248), .COUT(n27249));
    defparam sub_2057_add_2_5.INIT0 = 16'h5999;
    defparam sub_2057_add_2_5.INIT1 = 16'h5999;
    defparam sub_2057_add_2_5.INJECT1_0 = "NO";
    defparam sub_2057_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27247), .COUT(n27248));
    defparam sub_2057_add_2_3.INIT0 = 16'h5999;
    defparam sub_2057_add_2_3.INIT1 = 16'h5999;
    defparam sub_2057_add_2_3.INJECT1_0 = "NO";
    defparam sub_2057_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2057_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27247));
    defparam sub_2057_add_2_1.INIT0 = 16'h0000;
    defparam sub_2057_add_2_1.INIT1 = 16'h5999;
    defparam sub_2057_add_2_1.INJECT1_0 = "NO";
    defparam sub_2057_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27246), .S1(n8100));
    defparam sub_2059_add_2_33.INIT0 = 16'h5999;
    defparam sub_2059_add_2_33.INIT1 = 16'h0000;
    defparam sub_2059_add_2_33.INJECT1_0 = "NO";
    defparam sub_2059_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27245), .COUT(n27246));
    defparam sub_2059_add_2_31.INIT0 = 16'h5999;
    defparam sub_2059_add_2_31.INIT1 = 16'h5999;
    defparam sub_2059_add_2_31.INJECT1_0 = "NO";
    defparam sub_2059_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27244), .COUT(n27245));
    defparam sub_2059_add_2_29.INIT0 = 16'h5999;
    defparam sub_2059_add_2_29.INIT1 = 16'h5999;
    defparam sub_2059_add_2_29.INJECT1_0 = "NO";
    defparam sub_2059_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27243), .COUT(n27244));
    defparam sub_2059_add_2_27.INIT0 = 16'h5999;
    defparam sub_2059_add_2_27.INIT1 = 16'h5999;
    defparam sub_2059_add_2_27.INJECT1_0 = "NO";
    defparam sub_2059_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27242), .COUT(n27243));
    defparam sub_2059_add_2_25.INIT0 = 16'h5999;
    defparam sub_2059_add_2_25.INIT1 = 16'h5999;
    defparam sub_2059_add_2_25.INJECT1_0 = "NO";
    defparam sub_2059_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27241), .COUT(n27242));
    defparam sub_2059_add_2_23.INIT0 = 16'h5999;
    defparam sub_2059_add_2_23.INIT1 = 16'h5999;
    defparam sub_2059_add_2_23.INJECT1_0 = "NO";
    defparam sub_2059_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27240), .COUT(n27241));
    defparam sub_2059_add_2_21.INIT0 = 16'h5999;
    defparam sub_2059_add_2_21.INIT1 = 16'h5999;
    defparam sub_2059_add_2_21.INJECT1_0 = "NO";
    defparam sub_2059_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27239), .COUT(n27240));
    defparam sub_2059_add_2_19.INIT0 = 16'h5999;
    defparam sub_2059_add_2_19.INIT1 = 16'h5999;
    defparam sub_2059_add_2_19.INJECT1_0 = "NO";
    defparam sub_2059_add_2_19.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n32130), .CD(n16775), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_2059_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27238), .COUT(n27239));
    defparam sub_2059_add_2_17.INIT0 = 16'h5999;
    defparam sub_2059_add_2_17.INIT1 = 16'h5999;
    defparam sub_2059_add_2_17.INJECT1_0 = "NO";
    defparam sub_2059_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27237), .COUT(n27238));
    defparam sub_2059_add_2_15.INIT0 = 16'h5999;
    defparam sub_2059_add_2_15.INIT1 = 16'h5999;
    defparam sub_2059_add_2_15.INJECT1_0 = "NO";
    defparam sub_2059_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27236), .COUT(n27237));
    defparam sub_2059_add_2_13.INIT0 = 16'h5999;
    defparam sub_2059_add_2_13.INIT1 = 16'h5999;
    defparam sub_2059_add_2_13.INJECT1_0 = "NO";
    defparam sub_2059_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27235), .COUT(n27236));
    defparam sub_2059_add_2_11.INIT0 = 16'h5999;
    defparam sub_2059_add_2_11.INIT1 = 16'h5999;
    defparam sub_2059_add_2_11.INJECT1_0 = "NO";
    defparam sub_2059_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27234), .COUT(n27235));
    defparam sub_2059_add_2_9.INIT0 = 16'h5999;
    defparam sub_2059_add_2_9.INIT1 = 16'h5999;
    defparam sub_2059_add_2_9.INJECT1_0 = "NO";
    defparam sub_2059_add_2_9.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27694), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_33.INIT1 = 16'h0000;
    defparam count_2663_add_4_33.INJECT1_0 = "NO";
    defparam count_2663_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27693), .COUT(n27694), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2663_add_4_31.INJECT1_0 = "NO";
    defparam count_2663_add_4_31.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27233), .COUT(n27234));
    defparam sub_2059_add_2_7.INIT0 = 16'h5999;
    defparam sub_2059_add_2_7.INIT1 = 16'h5999;
    defparam sub_2059_add_2_7.INJECT1_0 = "NO";
    defparam sub_2059_add_2_7.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27692), .COUT(n27693), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2663_add_4_29.INJECT1_0 = "NO";
    defparam count_2663_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27691), .COUT(n27692), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2663_add_4_27.INJECT1_0 = "NO";
    defparam count_2663_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27690), .COUT(n27691), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2663_add_4_25.INJECT1_0 = "NO";
    defparam count_2663_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27232), .COUT(n27233));
    defparam sub_2059_add_2_5.INIT0 = 16'h5999;
    defparam sub_2059_add_2_5.INIT1 = 16'h5999;
    defparam sub_2059_add_2_5.INJECT1_0 = "NO";
    defparam sub_2059_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2059_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27231), .COUT(n27232));
    defparam sub_2059_add_2_3.INIT0 = 16'h5999;
    defparam sub_2059_add_2_3.INIT1 = 16'h5999;
    defparam sub_2059_add_2_3.INJECT1_0 = "NO";
    defparam sub_2059_add_2_3.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27689), .COUT(n27690), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2663_add_4_23.INJECT1_0 = "NO";
    defparam count_2663_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27688), .COUT(n27689), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2663_add_4_21.INJECT1_0 = "NO";
    defparam count_2663_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27687), .COUT(n27688), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2663_add_4_19.INJECT1_0 = "NO";
    defparam count_2663_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27686), .COUT(n27687), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2663_add_4_17.INJECT1_0 = "NO";
    defparam count_2663_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27685), .COUT(n27686), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2663_add_4_15.INJECT1_0 = "NO";
    defparam count_2663_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27684), .COUT(n27685), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2663_add_4_13.INJECT1_0 = "NO";
    defparam count_2663_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27683), .COUT(n27684), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2663_add_4_11.INJECT1_0 = "NO";
    defparam count_2663_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27682), .COUT(n27683), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2663_add_4_9.INJECT1_0 = "NO";
    defparam count_2663_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27681), .COUT(n27682), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2663_add_4_7.INJECT1_0 = "NO";
    defparam count_2663_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27680), .COUT(n27681), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2663_add_4_5.INJECT1_0 = "NO";
    defparam count_2663_add_4_5.INJECT1_1 = "NO";
    FD1S3IX count_2663__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i1.GSR = "ENABLED";
    CCU2D count_2663_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27679), .COUT(n27680), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2663_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2663_add_4_3.INJECT1_0 = "NO";
    defparam count_2663_add_4_3.INJECT1_1 = "NO";
    FD1S3IX count_2663__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i2.GSR = "ENABLED";
    FD1S3IX count_2663__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i3.GSR = "ENABLED";
    FD1S3IX count_2663__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i4.GSR = "ENABLED";
    FD1S3IX count_2663__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i5.GSR = "ENABLED";
    FD1S3IX count_2663__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i6.GSR = "ENABLED";
    FD1S3IX count_2663__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i7.GSR = "ENABLED";
    FD1S3IX count_2663__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i8.GSR = "ENABLED";
    FD1S3IX count_2663__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i9.GSR = "ENABLED";
    FD1S3IX count_2663__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i10.GSR = "ENABLED";
    FD1S3IX count_2663__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i11.GSR = "ENABLED";
    FD1S3IX count_2663__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i12.GSR = "ENABLED";
    FD1S3IX count_2663__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i13.GSR = "ENABLED";
    FD1S3IX count_2663__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i14.GSR = "ENABLED";
    FD1S3IX count_2663__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i15.GSR = "ENABLED";
    FD1S3IX count_2663__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i16.GSR = "ENABLED";
    FD1S3IX count_2663__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i17.GSR = "ENABLED";
    FD1S3IX count_2663__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i18.GSR = "ENABLED";
    FD1S3IX count_2663__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i19.GSR = "ENABLED";
    FD1S3IX count_2663__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i20.GSR = "ENABLED";
    FD1S3IX count_2663__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i21.GSR = "ENABLED";
    FD1S3IX count_2663__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i22.GSR = "ENABLED";
    FD1S3IX count_2663__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i23.GSR = "ENABLED";
    FD1S3IX count_2663__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i24.GSR = "ENABLED";
    FD1S3IX count_2663__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i25.GSR = "ENABLED";
    FD1S3IX count_2663__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i26.GSR = "ENABLED";
    FD1S3IX count_2663__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i27.GSR = "ENABLED";
    FD1S3IX count_2663__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i28.GSR = "ENABLED";
    FD1S3IX count_2663__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i29.GSR = "ENABLED";
    FD1S3IX count_2663__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i30.GSR = "ENABLED";
    FD1S3IX count_2663__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n32130), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663__i31.GSR = "ENABLED";
    CCU2D sub_2059_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27231));
    defparam sub_2059_add_2_1.INIT0 = 16'h0000;
    defparam sub_2059_add_2_1.INIT1 = 16'h5999;
    defparam sub_2059_add_2_1.INJECT1_0 = "NO";
    defparam sub_2059_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2663_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27679), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2663_add_4_1.INIT0 = 16'hF000;
    defparam count_2663_add_4_1.INIT1 = 16'h0555;
    defparam count_2663_add_4_1.INJECT1_0 = "NO";
    defparam count_2663_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_2060_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27230), .S1(n8134));
    defparam sub_2060_add_2_33.INIT0 = 16'hf555;
    defparam sub_2060_add_2_33.INIT1 = 16'h0000;
    defparam sub_2060_add_2_33.INJECT1_0 = "NO";
    defparam sub_2060_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2060_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27229), .COUT(n27230));
    defparam sub_2060_add_2_31.INIT0 = 16'hf555;
    defparam sub_2060_add_2_31.INIT1 = 16'hf555;
    defparam sub_2060_add_2_31.INJECT1_0 = "NO";
    defparam sub_2060_add_2_31.INJECT1_1 = "NO";
    LUT4 i1024_2_lut_rep_309 (.A(n8100), .B(n34065), .Z(n32130)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i1024_2_lut_rep_309.init = 16'heeee;
    LUT4 i10083_2_lut_3_lut (.A(n8100), .B(n34065), .C(n8134), .Z(n16775)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i10083_2_lut_3_lut.init = 16'he0e0;
    CCU2D sub_2060_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27228), .COUT(n27229));
    defparam sub_2060_add_2_29.INIT0 = 16'hf555;
    defparam sub_2060_add_2_29.INIT1 = 16'hf555;
    defparam sub_2060_add_2_29.INJECT1_0 = "NO";
    defparam sub_2060_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2060_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27227), .COUT(n27228));
    defparam sub_2060_add_2_27.INIT0 = 16'hf555;
    defparam sub_2060_add_2_27.INIT1 = 16'hf555;
    defparam sub_2060_add_2_27.INJECT1_0 = "NO";
    defparam sub_2060_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2060_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27226), .COUT(n27227));
    defparam sub_2060_add_2_25.INIT0 = 16'hf555;
    defparam sub_2060_add_2_25.INIT1 = 16'hf555;
    defparam sub_2060_add_2_25.INJECT1_0 = "NO";
    defparam sub_2060_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2060_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27225), .COUT(n27226));
    defparam sub_2060_add_2_23.INIT0 = 16'hf555;
    defparam sub_2060_add_2_23.INIT1 = 16'hf555;
    defparam sub_2060_add_2_23.INJECT1_0 = "NO";
    defparam sub_2060_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2060_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27224), .COUT(n27225));
    defparam sub_2060_add_2_21.INIT0 = 16'hf555;
    defparam sub_2060_add_2_21.INIT1 = 16'hf555;
    defparam sub_2060_add_2_21.INJECT1_0 = "NO";
    defparam sub_2060_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2060_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27223), .COUT(n27224));
    defparam sub_2060_add_2_19.INIT0 = 16'hf555;
    defparam sub_2060_add_2_19.INIT1 = 16'hf555;
    defparam sub_2060_add_2_19.INJECT1_0 = "NO";
    defparam sub_2060_add_2_19.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module RCPeripheral
//

module RCPeripheral (n2, databus, \register_addr[0] , \read_value[25] , 
            n8, n32141, n2_adj_58, databus_out, n34064, read_value, 
            \read_value[9]_adj_60 , n52, n32164, \select[7] , n176, 
            n2_adj_61, n2_adj_62, \read_value[11]_adj_63 , n8_adj_64, 
            read_value_adj_287, read_value_adj_288, n46, n52_adj_129, 
            \read_value[21]_adj_130 , n8_adj_131, n2_adj_132, \read_value[20]_adj_133 , 
            n8_adj_134, \read_value[11]_adj_135 , rw, \read_value[20]_adj_136 , 
            read_size, \select[1] , n32284, \sendcount[1] , n12746, 
            n2_adj_137, \read_value[19]_adj_138 , n8_adj_139, \register_addr[1] , 
            \read_value[19]_adj_140 , n2_adj_141, \read_value[10]_adj_142 , 
            n8_adj_143, n3, n2_adj_144, \read_value[18]_adj_145 , n8_adj_146, 
            read_value_adj_289, n64, n19559, read_value_adj_290, n2_adj_163, 
            \read_value[18]_adj_164 , \read_value[3]_adj_165 , \read_value[3]_adj_166 , 
            n32161, n2_adj_167, \read_value[8]_adj_168 , n8_adj_169, 
            n3_adj_170, n2_adj_171, \read_value[17]_adj_172 , n8_adj_173, 
            \read_value[28]_adj_174 , n8_adj_175, \read_value[10]_adj_176 , 
            \read_value[17]_adj_177 , \register_addr[2] , \register_addr[5] , 
            n2_adj_178, \read_value[16]_adj_179 , n8_adj_180, \read_value[16]_adj_181 , 
            \read_value[13]_adj_182 , \read_value[8]_adj_183 , n2_adj_184, 
            \read_value[15]_adj_185 , n8_adj_186, \read_value[15]_adj_187 , 
            n32282, \read_size[2]_adj_188 , \register_addr[4] , \read_size[2]_adj_189 , 
            n2_adj_190, \read_value[2]_adj_191 , \read_value[2]_adj_192 , 
            \read_size[2]_adj_193 , \read_size[2]_adj_194 , n2_adj_195, 
            \read_value[14]_adj_196 , n8_adj_197, n3_adj_198, n10, \read_value[12]_adj_199 , 
            n8_adj_200, \read_value[1]_adj_201 , n3_adj_202, \read_value[1]_adj_203 , 
            \read_value[14]_adj_204 , n2_adj_205, \read_value[9]_adj_206 , 
            n8_adj_207, n2_adj_208, \read_value[13]_adj_209 , n8_adj_210, 
            \read_value[25]_adj_211 , \read_value[28]_adj_212 , n2_adj_213, 
            \read_value[27]_adj_214 , n8_adj_215, \read_value[27]_adj_216 , 
            \read_value[21]_adj_217 , n2_adj_218, \read_value[6]_adj_219 , 
            \read_value[6]_adj_220 , n2_adj_221, n32185, \read_value[24]_adj_222 , 
            n8_adj_223, n13, \read_size[0]_adj_224 , n9, n32215, n18, 
            \read_size[0]_adj_225 , \read_size[0]_adj_226 , n32182, \select[2] , 
            n14, \read_size[0]_adj_227 , n5, n32155, \read_size[0]_adj_228 , 
            \read_size[0]_adj_229 , \select[5] , n32203, n32178, \read_size[2]_adj_230 , 
            \reg_size[2] , n3_adj_231, \read_size[2]_adj_232 , n32251, 
            n2_adj_233, \read_value[26]_adj_234 , n8_adj_235, \read_value[26]_adj_236 , 
            \read_value[24]_adj_237 , \read_value[12]_adj_238 , n2_adj_239, 
            \read_value[0]_adj_240 , \read_value[0]_adj_241 , n3_adj_242, 
            n2_adj_243, \read_value[31]_adj_244 , n8_adj_245, \read_value[31]_adj_246 , 
            n2_adj_247, n2_adj_248, n2_adj_249, n29920, n2_adj_250, 
            \read_value[30]_adj_251 , n8_adj_252, \read_value[30]_adj_253 , 
            \read_value[7]_adj_254 , \read_value[7]_adj_255 , n2_adj_256, 
            \read_value[29]_adj_257 , n8_adj_258, \read_value[29]_adj_259 , 
            \read_value[4]_adj_260 , \read_value[4]_adj_261 , n2_adj_262, 
            \read_value[5]_adj_263 , \read_value[5]_adj_264 , \read_value[23]_adj_265 , 
            n8_adj_266, \read_value[23]_adj_267 , n3_adj_268, n3_adj_269, 
            n2_adj_270, \read_value[22]_adj_271 , n8_adj_272, \read_value[22]_adj_273 , 
            n2_adj_274, \count[6] , \count[5] , n29947, n5_adj_275, 
            GND_net, n30260, \count[8] , \count[9] , n30482, n32135, 
            n30304, n32302, \count[4] , n32245, n32301, n28333, 
            debug_c_c, rc_ch8_c, n32256, \count[1] , \count[2] , n32257, 
            \count[3] , n32218, n32258, n13605, \count[0] , n30001, 
            n29948, n28141, n28234, n32129, n32134, n30474, rc_ch7_c, 
            n30623, n28140, n32283, n28331, n32317, n13974, rc_ch4_c, 
            n28133, n30472, n28233, n32221, \count[9]_adj_276 , n32264, 
            n28330, n5_adj_277, \count[5]_adj_278 , n5_adj_279, \count[6]_adj_280 , 
            n32267, \count[8]_adj_281 , n13975, rc_ch3_c, n28132, 
            n28222, n32127, n30470, n30302, n28232, n32125, n32294, 
            \count[9]_adj_282 , \count[8]_adj_283 , \count[5]_adj_284 , 
            \count[6]_adj_285 , rc_ch2_c, n13976, n5_adj_286, n32293, 
            n41, n28329, n32296, n28144, n30308, n30465, n13977, 
            n30463, n32274, n28328, n32308, rc_ch1_c, n28231, n28129) /* synthesis syn_module_defined=1 */ ;
    input n2;
    output [31:0]databus;
    input \register_addr[0] ;
    input \read_value[25] ;
    input n8;
    input n32141;
    input n2_adj_58;
    input [31:0]databus_out;
    input n34064;
    input [31:0]read_value;
    input \read_value[9]_adj_60 ;
    input n52;
    input n32164;
    input \select[7] ;
    input n176;
    input n2_adj_61;
    input n2_adj_62;
    input \read_value[11]_adj_63 ;
    input n8_adj_64;
    input [31:0]read_value_adj_287;
    input [31:0]read_value_adj_288;
    input n46;
    input n52_adj_129;
    input \read_value[21]_adj_130 ;
    input n8_adj_131;
    input n2_adj_132;
    input \read_value[20]_adj_133 ;
    input n8_adj_134;
    input \read_value[11]_adj_135 ;
    input rw;
    input \read_value[20]_adj_136 ;
    input [2:0]read_size;
    input \select[1] ;
    output n32284;
    input \sendcount[1] ;
    output n12746;
    input n2_adj_137;
    input \read_value[19]_adj_138 ;
    input n8_adj_139;
    input \register_addr[1] ;
    input \read_value[19]_adj_140 ;
    input n2_adj_141;
    input \read_value[10]_adj_142 ;
    input n8_adj_143;
    input n3;
    input n2_adj_144;
    input \read_value[18]_adj_145 ;
    input n8_adj_146;
    input [7:0]read_value_adj_289;
    input n64;
    input n19559;
    input [7:0]read_value_adj_290;
    input n2_adj_163;
    input \read_value[18]_adj_164 ;
    input \read_value[3]_adj_165 ;
    input \read_value[3]_adj_166 ;
    input n32161;
    input n2_adj_167;
    input \read_value[8]_adj_168 ;
    input n8_adj_169;
    input n3_adj_170;
    input n2_adj_171;
    input \read_value[17]_adj_172 ;
    input n8_adj_173;
    input \read_value[28]_adj_174 ;
    input n8_adj_175;
    input \read_value[10]_adj_176 ;
    input \read_value[17]_adj_177 ;
    input \register_addr[2] ;
    input \register_addr[5] ;
    input n2_adj_178;
    input \read_value[16]_adj_179 ;
    input n8_adj_180;
    input \read_value[16]_adj_181 ;
    input \read_value[13]_adj_182 ;
    input \read_value[8]_adj_183 ;
    input n2_adj_184;
    input \read_value[15]_adj_185 ;
    input n8_adj_186;
    input \read_value[15]_adj_187 ;
    input n32282;
    input \read_size[2]_adj_188 ;
    input \register_addr[4] ;
    input \read_size[2]_adj_189 ;
    input n2_adj_190;
    input \read_value[2]_adj_191 ;
    input \read_value[2]_adj_192 ;
    input \read_size[2]_adj_193 ;
    input \read_size[2]_adj_194 ;
    input n2_adj_195;
    input \read_value[14]_adj_196 ;
    input n8_adj_197;
    input n3_adj_198;
    input n10;
    input \read_value[12]_adj_199 ;
    input n8_adj_200;
    input \read_value[1]_adj_201 ;
    input n3_adj_202;
    input \read_value[1]_adj_203 ;
    input \read_value[14]_adj_204 ;
    input n2_adj_205;
    input \read_value[9]_adj_206 ;
    input n8_adj_207;
    input n2_adj_208;
    input \read_value[13]_adj_209 ;
    input n8_adj_210;
    input \read_value[25]_adj_211 ;
    input \read_value[28]_adj_212 ;
    input n2_adj_213;
    input \read_value[27]_adj_214 ;
    input n8_adj_215;
    input \read_value[27]_adj_216 ;
    input \read_value[21]_adj_217 ;
    input n2_adj_218;
    input \read_value[6]_adj_219 ;
    input \read_value[6]_adj_220 ;
    input n2_adj_221;
    input n32185;
    input \read_value[24]_adj_222 ;
    input n8_adj_223;
    output n13;
    input \read_size[0]_adj_224 ;
    input n9;
    input n32215;
    output n18;
    input \read_size[0]_adj_225 ;
    input \read_size[0]_adj_226 ;
    input n32182;
    input \select[2] ;
    output n14;
    input \read_size[0]_adj_227 ;
    input n5;
    input n32155;
    input \read_size[0]_adj_228 ;
    input \read_size[0]_adj_229 ;
    input \select[5] ;
    input n32203;
    input n32178;
    input \read_size[2]_adj_230 ;
    output \reg_size[2] ;
    input n3_adj_231;
    input \read_size[2]_adj_232 ;
    input n32251;
    input n2_adj_233;
    input \read_value[26]_adj_234 ;
    input n8_adj_235;
    input \read_value[26]_adj_236 ;
    input \read_value[24]_adj_237 ;
    input \read_value[12]_adj_238 ;
    input n2_adj_239;
    input \read_value[0]_adj_240 ;
    input \read_value[0]_adj_241 ;
    input n3_adj_242;
    input n2_adj_243;
    input \read_value[31]_adj_244 ;
    input n8_adj_245;
    input \read_value[31]_adj_246 ;
    input n2_adj_247;
    input n2_adj_248;
    input n2_adj_249;
    output n29920;
    input n2_adj_250;
    input \read_value[30]_adj_251 ;
    input n8_adj_252;
    input \read_value[30]_adj_253 ;
    input \read_value[7]_adj_254 ;
    input \read_value[7]_adj_255 ;
    input n2_adj_256;
    input \read_value[29]_adj_257 ;
    input n8_adj_258;
    input \read_value[29]_adj_259 ;
    input \read_value[4]_adj_260 ;
    input \read_value[4]_adj_261 ;
    input n2_adj_262;
    input \read_value[5]_adj_263 ;
    input \read_value[5]_adj_264 ;
    input \read_value[23]_adj_265 ;
    input n8_adj_266;
    input \read_value[23]_adj_267 ;
    input n3_adj_268;
    input n3_adj_269;
    input n2_adj_270;
    input \read_value[22]_adj_271 ;
    input n8_adj_272;
    input \read_value[22]_adj_273 ;
    input n2_adj_274;
    output \count[6] ;
    output \count[5] ;
    output n29947;
    output n5_adj_275;
    input GND_net;
    output n30260;
    output \count[8] ;
    output \count[9] ;
    output n30482;
    input n32135;
    output n30304;
    input n32302;
    output \count[4] ;
    input n32245;
    output n32301;
    output n28333;
    input debug_c_c;
    input rc_ch8_c;
    output n32256;
    output \count[1] ;
    output \count[2] ;
    output n32257;
    output \count[3] ;
    output n32218;
    output n32258;
    input n13605;
    output \count[0] ;
    input n30001;
    input n29948;
    output n28141;
    input n28234;
    input n32129;
    input n32134;
    output n30474;
    input rc_ch7_c;
    output n30623;
    input n28140;
    output n32283;
    output n28331;
    output n32317;
    input n13974;
    input rc_ch4_c;
    output n28133;
    output n30472;
    input n28233;
    output n32221;
    output \count[9]_adj_276 ;
    output n32264;
    output n28330;
    output n5_adj_277;
    output \count[5]_adj_278 ;
    output n5_adj_279;
    output \count[6]_adj_280 ;
    output n32267;
    output \count[8]_adj_281 ;
    input n13975;
    input rc_ch3_c;
    output n28132;
    input n28222;
    input n32127;
    output n30470;
    output n30302;
    input n28232;
    input n32125;
    output n32294;
    output \count[9]_adj_282 ;
    output \count[8]_adj_283 ;
    output \count[5]_adj_284 ;
    output \count[6]_adj_285 ;
    input rc_ch2_c;
    input n13976;
    output n5_adj_286;
    output n32293;
    output n41;
    output n28329;
    output n32296;
    output n28144;
    output n30308;
    output n30465;
    input n13977;
    output n30463;
    output n32274;
    output n28328;
    output n32308;
    input rc_ch1_c;
    input n28231;
    output n28129;
    
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(455[15:21])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n13_c, n11, n5_c;
    wire [7:0]\register[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n31830;
    wire [7:0]\register[6] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n31829, n10_c, n13_adj_173, n11_adj_174, n5_adj_176, n5_adj_177, 
        n10_adj_179;
    wire [2:0]read_size_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(211[12:21])
    
    wire n31905, n13_adj_180, n11_adj_181, n31906;
    wire [7:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    wire [7:0]\register[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n31578, n13_adj_183, n11_adj_184, n5_adj_186;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(207[13:21])
    
    wire n31579, n10_adj_187, n10_adj_192, n13_adj_194, n13_adj_195, 
        n11_adj_196, n5_adj_198, n10_adj_199, n31908, n1105, n31909, 
        n31707, n13_adj_207, n11_adj_208, n5_adj_210, n10_adj_211, 
        n31576, n31575, n31577, n13_adj_217, n11_adj_218, n5_adj_220, 
        n5_adj_221, n10_adj_222, n31977, n1180, n31978, n7, n14_c, 
        n18_c, n13_adj_226, n11_adj_227, n5_adj_229, n10_adj_230, 
        n12, n15, n20, n7_adj_239;
    wire [7:0]read_value_adj_556;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(210[12:22])
    
    wire n18_adj_244, n12_adj_245, n46_adj_246, n31975, n13_adj_249, 
        n11_adj_250, n5_adj_252, n10_adj_253, n14_adj_256, n31974, 
        n31981, n31982, n31984, n1135, n31985, n13_adj_262, n11_adj_263, 
        n5_adj_265, n10_adj_266, n10_adj_270, n31526, n31523, n31527, 
        n26, n29998, n32, n13_adj_276, n11_adj_277, n5_adj_279_c, 
        n10_adj_280, n31706, n31709, n10_adj_287, n1120, n31710, 
        n32101, n32100, n31525, n31524, n32103, n32104, n13_adj_292, 
        n11_adj_293, n5_adj_295, n10_adj_296, n15_adj_305, n20_adj_306, 
        n7_adj_308, n18_adj_311, n12_adj_312, n13_adj_315, n11_adj_316, 
        n5_adj_318, n10_adj_319, n14_adj_324, n19, n8_adj_330, n18_adj_331, 
        n12_adj_332, n16, n10_adj_334, n14_adj_337, n13_adj_349, n11_adj_350, 
        n5_adj_352, n13_adj_355, n11_adj_356, n11_adj_368, n1150, 
        n31833, n31832, n32105, n32102, n32106, n5_adj_371, n31521, 
        n13_adj_372, n11_adj_373, n5_adj_375, n31522, n10_adj_376, 
        n1165, n31986, n31983, n31987, n15_adj_384, n20_adj_385, 
        n7_adj_387, n31979, n31976, n31980, n13_adj_389, n11_adj_390, 
        n5_adj_392, n31712, n31835, n31581, n18_adj_395, n12_adj_396, 
        n10_adj_397, n16_adj_402, n12_adj_408, n6, n1, n14_adj_414, 
        n13_adj_418, n11_adj_419, n5_adj_421, n10_adj_422, n31910, 
        n31907, n31911, n15_adj_436, n20_adj_437, n7_adj_439, n18_adj_442, 
        n12_adj_443, n14_adj_445, n31834, n31831, n13_adj_451, n11_adj_452, 
        n5_adj_454, n10_adj_455, n15_adj_461, n20_adj_462, n7_adj_464, 
        n13_adj_465, n11_adj_466, n5_adj_468, n15_adj_469, n20_adj_470, 
        n13_adj_474, n11_adj_475, n5_adj_477, n10_adj_478, n13_adj_486, 
        n11_adj_487, n5_adj_489, n10_adj_490, n31711, n31708, n18_adj_496, 
        n12_adj_497, n15_adj_500, n20_adj_501, n7_adj_503, n18_adj_506, 
        n12_adj_507, n10_adj_508, n14_adj_515, n14_adj_518, n13_adj_520, 
        n11_adj_521, n5_adj_523, n10_adj_528, n31580;
    
    LUT4 i7_4_lut (.A(n13_c), .B(n11), .C(n2), .D(n5_c), .Z(databus[25])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 register_addr_1__bdd_3_lut_23616 (.A(\register_addr[0] ), .B(\register[4] [3]), 
         .C(\register[5] [3]), .Z(n31830)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23616.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_23615 (.A(\register[6] [3]), .B(\register_addr[0] ), 
         .Z(n31829)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23615.init = 16'h2222;
    LUT4 i5_4_lut (.A(\read_value[25] ), .B(n10_c), .C(n8), .D(n32141), 
         .Z(n13_c)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut.init = 16'hfefc;
    LUT4 i7_4_lut_adj_318 (.A(n13_adj_173), .B(n11_adj_174), .C(n2_adj_58), 
         .D(n5_adj_176), .Z(databus[28])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_318.init = 16'hfffe;
    LUT4 Select_4266_i5_2_lut (.A(databus_out[12]), .B(n34064), .Z(n5_adj_177)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4266_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut (.A(read_value[9]), .B(\read_value[9]_adj_60 ), .C(n52), 
         .D(n32164), .Z(n10_adj_179)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut.init = 16'heca0;
    FD1S3AX read_size_i1 (.D(n176), .CK(\select[7] ), .Q(read_size_c[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_size_i1.GSR = "ENABLED";
    LUT4 register_addr_1__bdd_2_lut_23648 (.A(\register[6] [0]), .B(\register_addr[0] ), 
         .Z(n31905)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23648.init = 16'h2222;
    LUT4 i7_4_lut_adj_319 (.A(n13_adj_180), .B(n11_adj_181), .C(n2_adj_61), 
         .D(n5_adj_177), .Z(databus[12])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_319.init = 16'hfffe;
    LUT4 register_addr_1__bdd_3_lut_23649 (.A(\register_addr[0] ), .B(\register[4] [0]), 
         .C(\register[5] [0]), .Z(n31906)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23649.init = 16'he4e4;
    LUT4 \register_1[[4__bdd_3_lut_23731  (.A(\register[2] [4]), .B(\register[3] [4]), 
         .C(\register_addr[0] ), .Z(n31578)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[4__bdd_3_lut_23731 .init = 16'hcaca;
    LUT4 i7_4_lut_adj_320 (.A(n13_adj_183), .B(n11_adj_184), .C(n2_adj_62), 
         .D(n5_adj_186), .Z(databus[11])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_320.init = 16'hfffe;
    LUT4 \register_1[[4__bdd_2_lut_23732  (.A(\register[1] [4]), .B(\register_addr[0] ), 
         .Z(n31579)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[4__bdd_2_lut_23732 .init = 16'h8888;
    LUT4 i5_4_lut_adj_321 (.A(\read_value[11]_adj_63 ), .B(n10_adj_187), 
         .C(n8_adj_64), .D(n32141), .Z(n13_adj_183)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_321.init = 16'hfefc;
    LUT4 i3_4_lut (.A(read_value_adj_287[11]), .B(read_value_adj_288[11]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_184)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut.init = 16'heca0;
    LUT4 i5_4_lut_adj_322 (.A(\read_value[21]_adj_130 ), .B(n10_adj_192), 
         .C(n8_adj_131), .D(n32141), .Z(n13_adj_194)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_322.init = 16'hfefc;
    LUT4 i7_4_lut_adj_323 (.A(n13_adj_195), .B(n11_adj_196), .C(n2_adj_132), 
         .D(n5_adj_198), .Z(databus[20])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_323.init = 16'hfffe;
    LUT4 i5_4_lut_adj_324 (.A(\read_value[20]_adj_133 ), .B(n10_adj_199), 
         .C(n8_adj_134), .D(n32141), .Z(n13_adj_195)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_324.init = 16'hfefc;
    LUT4 Select_4269_i5_2_lut (.A(databus_out[11]), .B(n34064), .Z(n5_adj_186)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4269_i5_2_lut.init = 16'h2222;
    LUT4 i3_4_lut_adj_325 (.A(read_value_adj_287[20]), .B(read_value_adj_288[20]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_196)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_325.init = 16'heca0;
    LUT4 i2_4_lut_adj_326 (.A(read_value[11]), .B(\read_value[11]_adj_135 ), 
         .C(n52), .D(n32164), .Z(n10_adj_187)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_326.init = 16'heca0;
    LUT4 n1105_bdd_3_lut_23627 (.A(\register[2] [0]), .B(\register[3] [0]), 
         .C(\register_addr[0] ), .Z(n31908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1105_bdd_3_lut_23627.init = 16'hcaca;
    LUT4 n1105_bdd_3_lut_23634 (.A(n1105), .B(\register_addr[0] ), .C(\register[1] [0]), 
         .Z(n31909)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1105_bdd_3_lut_23634.init = 16'he2e2;
    LUT4 Select_4242_i5_2_lut (.A(databus_out[20]), .B(rw), .Z(n5_adj_198)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4242_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_327 (.A(read_value[20]), .B(\read_value[20]_adj_136 ), 
         .C(n52), .D(n32164), .Z(n10_adj_199)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_327.init = 16'heca0;
    LUT4 Select_4296_i1_2_lut_rep_463 (.A(read_size[1]), .B(\select[1] ), 
         .Z(n32284)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4296_i1_2_lut_rep_463.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(read_size[1]), .B(\select[1] ), .C(\sendcount[1] ), 
         .Z(n12746)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7878;
    LUT4 register_addr_1__bdd_3_lut_23598 (.A(\register_addr[0] ), .B(\register[4] [1]), 
         .C(\register[5] [1]), .Z(n31707)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23598.init = 16'he4e4;
    LUT4 i7_4_lut_adj_328 (.A(n13_adj_207), .B(n11_adj_208), .C(n2_adj_137), 
         .D(n5_adj_210), .Z(databus[19])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_328.init = 16'hfffe;
    LUT4 i5_4_lut_adj_329 (.A(\read_value[19]_adj_138 ), .B(n10_adj_211), 
         .C(n8_adj_139), .D(n32141), .Z(n13_adj_207)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_329.init = 16'hfefc;
    LUT4 i3_4_lut_adj_330 (.A(read_value_adj_287[19]), .B(read_value_adj_288[19]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_208)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_330.init = 16'heca0;
    PFUMX i23455 (.BLUT(n31576), .ALUT(n31575), .C0(\register_addr[1] ), 
          .Z(n31577));
    LUT4 Select_4245_i5_2_lut (.A(databus_out[19]), .B(rw), .Z(n5_adj_210)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4245_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_331 (.A(read_value[19]), .B(\read_value[19]_adj_140 ), 
         .C(n52), .D(n32164), .Z(n10_adj_211)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_331.init = 16'heca0;
    LUT4 i7_4_lut_adj_332 (.A(n13_adj_217), .B(n11_adj_218), .C(n2_adj_141), 
         .D(n5_adj_220), .Z(databus[10])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_332.init = 16'hfffe;
    LUT4 Select_4263_i5_2_lut (.A(databus_out[13]), .B(rw), .Z(n5_adj_221)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4263_i5_2_lut.init = 16'h2222;
    LUT4 i5_4_lut_adj_333 (.A(\read_value[10]_adj_142 ), .B(n10_adj_222), 
         .C(n8_adj_143), .D(n32141), .Z(n13_adj_217)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_333.init = 16'hfefc;
    LUT4 i3_4_lut_adj_334 (.A(read_value_adj_287[10]), .B(read_value_adj_288[10]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_218)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_334.init = 16'heca0;
    LUT4 n1180_bdd_3_lut_23658 (.A(\register[2] [7]), .B(\register[3] [7]), 
         .C(\register_addr[0] ), .Z(n31977)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1180_bdd_3_lut_23658.init = 16'hcaca;
    LUT4 n1180_bdd_3_lut_24275 (.A(n1180), .B(\register_addr[0] ), .C(\register[1] [7]), 
         .Z(n31978)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1180_bdd_3_lut_24275.init = 16'he2e2;
    LUT4 Select_4282_i7_2_lut (.A(databus_out[4]), .B(n34064), .Z(n7)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4282_i7_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_335 (.A(read_value_adj_287[4]), .B(n14_c), .C(n3), 
         .D(n46), .Z(n18_c)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_335.init = 16'hfefc;
    LUT4 i7_4_lut_adj_336 (.A(n13_adj_226), .B(n11_adj_227), .C(n2_adj_144), 
         .D(n5_adj_229), .Z(databus[18])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_336.init = 16'hfffe;
    LUT4 i5_4_lut_adj_337 (.A(\read_value[18]_adj_145 ), .B(n10_adj_230), 
         .C(n8_adj_146), .D(n32141), .Z(n13_adj_226)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_337.init = 16'hfefc;
    LUT4 i3_4_lut_adj_338 (.A(read_value_adj_287[18]), .B(read_value_adj_288[18]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_227)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_338.init = 16'heca0;
    LUT4 i1_4_lut (.A(read_value_adj_288[4]), .B(read_value_adj_289[4]), 
         .C(n52_adj_129), .D(n64), .Z(n12)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i3_4_lut_adj_339 (.A(read_value[4]), .B(n19559), .C(n52), .D(read_value_adj_290[4]), 
         .Z(n14_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_339.init = 16'heca0;
    LUT4 Select_4248_i5_2_lut (.A(databus_out[18]), .B(rw), .Z(n5_adj_229)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4248_i5_2_lut.init = 16'h2222;
    LUT4 i10_4_lut (.A(n15), .B(n20), .C(n2_adj_163), .D(n7_adj_239), 
         .Z(databus[3])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_340 (.A(read_value[18]), .B(\read_value[18]_adj_164 ), 
         .C(n52), .D(n32164), .Z(n10_adj_230)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_340.init = 16'heca0;
    LUT4 i4_4_lut (.A(\read_value[3]_adj_165 ), .B(\read_value[3]_adj_166 ), 
         .C(n32164), .D(n32161), .Z(n15)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut.init = 16'heca0;
    LUT4 i9_4_lut (.A(read_value_adj_556[3]), .B(n18_adj_244), .C(n12_adj_245), 
         .D(n46_adj_246), .Z(n20)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut.init = 16'hfefc;
    LUT4 register_addr_1__bdd_3_lut_23664 (.A(\register_addr[0] ), .B(\register[4] [7]), 
         .C(\register[5] [7]), .Z(n31975)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23664.init = 16'he4e4;
    LUT4 i3_4_lut_adj_341 (.A(read_value_adj_287[25]), .B(read_value_adj_288[25]), 
         .C(n46), .D(n52_adj_129), .Z(n11)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_341.init = 16'heca0;
    LUT4 i7_4_lut_adj_342 (.A(n13_adj_249), .B(n11_adj_250), .C(n2_adj_167), 
         .D(n5_adj_252), .Z(databus[8])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_342.init = 16'hfffe;
    LUT4 Select_4283_i7_2_lut (.A(databus_out[3]), .B(n34064), .Z(n7_adj_239)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4283_i7_2_lut.init = 16'h2222;
    LUT4 Select_4272_i5_2_lut (.A(databus_out[10]), .B(rw), .Z(n5_adj_220)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4272_i5_2_lut.init = 16'h2222;
    LUT4 i5_4_lut_adj_343 (.A(\read_value[8]_adj_168 ), .B(n10_adj_253), 
         .C(n8_adj_169), .D(n32141), .Z(n13_adj_249)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_343.init = 16'hfefc;
    LUT4 i7_4_lut_adj_344 (.A(read_value_adj_287[3]), .B(n14_adj_256), .C(n3_adj_170), 
         .D(n46), .Z(n18_adj_244)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_344.init = 16'hfefc;
    LUT4 i1_4_lut_adj_345 (.A(read_value_adj_288[3]), .B(read_value_adj_289[3]), 
         .C(n52_adj_129), .D(n64), .Z(n12_adj_245)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_345.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_23663 (.A(\register[6] [7]), .B(\register_addr[0] ), 
         .Z(n31974)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23663.init = 16'h2222;
    LUT4 i3_4_lut_adj_346 (.A(read_value[3]), .B(n19559), .C(n52), .D(read_value_adj_290[3]), 
         .Z(n14_adj_256)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_346.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_23715 (.A(\register[6] [2]), .B(\register_addr[0] ), 
         .Z(n31981)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23715.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut_23716 (.A(\register_addr[0] ), .B(\register[4] [2]), 
         .C(\register[5] [2]), .Z(n31982)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23716.init = 16'he4e4;
    LUT4 n1135_bdd_3_lut_23667 (.A(\register[2] [2]), .B(\register[3] [2]), 
         .C(\register_addr[0] ), .Z(n31984)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1135_bdd_3_lut_23667.init = 16'hcaca;
    LUT4 n1135_bdd_3_lut_24269 (.A(n1135), .B(\register_addr[0] ), .C(\register[1] [2]), 
         .Z(n31985)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1135_bdd_3_lut_24269.init = 16'he2e2;
    LUT4 i7_4_lut_adj_347 (.A(n13_adj_262), .B(n11_adj_263), .C(n2_adj_171), 
         .D(n5_adj_265), .Z(databus[17])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_347.init = 16'hfffe;
    LUT4 i5_4_lut_adj_348 (.A(\read_value[17]_adj_172 ), .B(n10_adj_266), 
         .C(n8_adj_173), .D(n32141), .Z(n13_adj_262)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_348.init = 16'hfefc;
    LUT4 i3_4_lut_adj_349 (.A(read_value_adj_287[17]), .B(read_value_adj_288[17]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_263)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_349.init = 16'heca0;
    LUT4 i5_4_lut_adj_350 (.A(\read_value[28]_adj_174 ), .B(n10_adj_270), 
         .C(n8_adj_175), .D(n32141), .Z(n13_adj_173)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_350.init = 16'hfefc;
    LUT4 i2_4_lut_adj_351 (.A(read_value[10]), .B(\read_value[10]_adj_176 ), 
         .C(n52), .D(n32164), .Z(n10_adj_222)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_351.init = 16'heca0;
    LUT4 Select_4251_i5_2_lut (.A(databus_out[17]), .B(rw), .Z(n5_adj_265)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4251_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_352 (.A(read_value[17]), .B(\read_value[17]_adj_177 ), 
         .C(n52), .D(n32164), .Z(n10_adj_266)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_352.init = 16'heca0;
    L6MUX21 i23418 (.D0(n31526), .D1(n31523), .SD(\register_addr[2] ), 
            .Z(n31527));
    PFUMX i45 (.BLUT(n26), .ALUT(n29998), .C0(\register_addr[5] ), .Z(n32));
    LUT4 i7_4_lut_adj_353 (.A(n13_adj_276), .B(n11_adj_277), .C(n2_adj_178), 
         .D(n5_adj_279_c), .Z(databus[16])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_353.init = 16'hfffe;
    LUT4 i5_4_lut_adj_354 (.A(\read_value[16]_adj_179 ), .B(n10_adj_280), 
         .C(n8_adj_180), .D(n32141), .Z(n13_adj_276)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_354.init = 16'hfefc;
    LUT4 i3_4_lut_adj_355 (.A(read_value_adj_287[16]), .B(read_value_adj_288[16]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_277)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_355.init = 16'heca0;
    LUT4 Select_4254_i5_2_lut (.A(databus_out[16]), .B(rw), .Z(n5_adj_279_c)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4254_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_356 (.A(read_value[16]), .B(\read_value[16]_adj_181 ), 
         .C(n52), .D(n32164), .Z(n10_adj_280)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_356.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_23597 (.A(\register[6] [1]), .B(\register_addr[0] ), 
         .Z(n31706)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23597.init = 16'h2222;
    LUT4 n1120_bdd_3_lut_23537 (.A(\register[2] [1]), .B(\register[3] [1]), 
         .C(\register_addr[0] ), .Z(n31709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1120_bdd_3_lut_23537.init = 16'hcaca;
    LUT4 i2_4_lut_adj_357 (.A(read_value[13]), .B(\read_value[13]_adj_182 ), 
         .C(n52), .D(n32164), .Z(n10_adj_287)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_357.init = 16'heca0;
    LUT4 n1120_bdd_3_lut_23702 (.A(n1120), .B(\register_addr[0] ), .C(\register[1] [1]), 
         .Z(n31710)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1120_bdd_3_lut_23702.init = 16'he2e2;
    LUT4 i3_4_lut_adj_358 (.A(read_value_adj_287[8]), .B(read_value_adj_288[8]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_250)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_358.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut (.A(\register_addr[0] ), .B(\register[4] [5]), 
         .C(\register[5] [5]), .Z(n32101)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut.init = 16'he4e4;
    LUT4 Select_4278_i5_2_lut (.A(databus_out[8]), .B(rw), .Z(n5_adj_252)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4278_i5_2_lut.init = 16'h2222;
    LUT4 register_addr_1__bdd_2_lut (.A(\register[6] [5]), .B(\register_addr[0] ), 
         .Z(n32100)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut.init = 16'h2222;
    PFUMX i23416 (.BLUT(n31525), .ALUT(n31524), .C0(\register_addr[1] ), 
          .Z(n31526));
    LUT4 \register_1[[5__bdd_3_lut_24244  (.A(\register[2] [5]), .B(\register[3] [5]), 
         .C(\register_addr[0] ), .Z(n32103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[5__bdd_3_lut_24244 .init = 16'hcaca;
    LUT4 i2_4_lut_adj_359 (.A(read_value[8]), .B(\read_value[8]_adj_183 ), 
         .C(n52), .D(n32164), .Z(n10_adj_253)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_359.init = 16'heca0;
    LUT4 \register_1[[5__bdd_2_lut_24245  (.A(\register[1] [5]), .B(\register_addr[0] ), 
         .Z(n32104)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[5__bdd_2_lut_24245 .init = 16'h8888;
    LUT4 n1165_bdd_3_lut_23415 (.A(\register[2] [6]), .B(\register[3] [6]), 
         .C(\register_addr[0] ), .Z(n31524)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1165_bdd_3_lut_23415.init = 16'hcaca;
    LUT4 i7_4_lut_adj_360 (.A(n13_adj_292), .B(n11_adj_293), .C(n2_adj_184), 
         .D(n5_adj_295), .Z(databus[15])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_360.init = 16'hfffe;
    LUT4 i5_4_lut_adj_361 (.A(\read_value[15]_adj_185 ), .B(n10_adj_296), 
         .C(n8_adj_186), .D(n32141), .Z(n13_adj_292)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_361.init = 16'hfefc;
    LUT4 i3_4_lut_adj_362 (.A(read_value_adj_287[15]), .B(read_value_adj_288[15]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_293)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_362.init = 16'heca0;
    LUT4 i3_4_lut_adj_363 (.A(read_value_adj_287[28]), .B(read_value_adj_288[28]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_174)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_363.init = 16'heca0;
    LUT4 Select_4257_i5_2_lut (.A(databus_out[15]), .B(rw), .Z(n5_adj_295)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4257_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_364 (.A(read_value[15]), .B(\read_value[15]_adj_187 ), 
         .C(n52), .D(n32164), .Z(n10_adj_296)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_364.init = 16'heca0;
    LUT4 i47_4_lut (.A(n32282), .B(\read_size[2]_adj_188 ), .C(\register_addr[4] ), 
         .D(\read_size[2]_adj_189 ), .Z(n26)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i47_4_lut.init = 16'h4540;
    LUT4 i10_4_lut_adj_365 (.A(n15_adj_305), .B(n20_adj_306), .C(n2_adj_190), 
         .D(n7_adj_308), .Z(databus[2])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_365.init = 16'hfffe;
    LUT4 i4_4_lut_adj_366 (.A(\read_value[2]_adj_191 ), .B(\read_value[2]_adj_192 ), 
         .C(n32164), .D(n32161), .Z(n15_adj_305)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_366.init = 16'heca0;
    LUT4 i9_4_lut_adj_367 (.A(read_value_adj_556[2]), .B(n18_adj_311), .C(n12_adj_312), 
         .D(n46_adj_246), .Z(n20_adj_306)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_367.init = 16'hfefc;
    LUT4 i1_4_lut_adj_368 (.A(\read_size[2]_adj_193 ), .B(n32282), .C(\read_size[2]_adj_194 ), 
         .D(\register_addr[4] ), .Z(n29998)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_368.init = 16'h3022;
    LUT4 i7_4_lut_adj_369 (.A(n13_adj_315), .B(n11_adj_316), .C(n2_adj_195), 
         .D(n5_adj_318), .Z(databus[14])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_369.init = 16'hfffe;
    LUT4 Select_4284_i7_2_lut (.A(databus_out[2]), .B(n34064), .Z(n7_adj_308)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4284_i7_2_lut.init = 16'h2222;
    LUT4 i5_4_lut_adj_370 (.A(\read_value[14]_adj_196 ), .B(n10_adj_319), 
         .C(n8_adj_197), .D(n32141), .Z(n13_adj_315)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_370.init = 16'hfefc;
    LUT4 i3_4_lut_adj_371 (.A(read_value_adj_287[14]), .B(read_value_adj_288[14]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_316)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_371.init = 16'heca0;
    LUT4 i7_4_lut_adj_372 (.A(read_value_adj_287[2]), .B(n14_adj_324), .C(n3_adj_198), 
         .D(n46), .Z(n18_adj_311)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_372.init = 16'hfefc;
    LUT4 i1_4_lut_adj_373 (.A(read_value_adj_288[2]), .B(read_value_adj_289[2]), 
         .C(n52_adj_129), .D(n64), .Z(n12_adj_312)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_373.init = 16'heca0;
    LUT4 i3_4_lut_adj_374 (.A(read_value[2]), .B(n19559), .C(n52), .D(read_value_adj_290[2]), 
         .Z(n14_adj_324)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_374.init = 16'heca0;
    LUT4 i10_4_lut_adj_375 (.A(n19), .B(n8_adj_330), .C(n18_adj_331), 
         .D(n12_adj_332), .Z(databus[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_375.init = 16'hfffe;
    LUT4 i8_4_lut (.A(read_value_adj_556[1]), .B(n16), .C(n10), .D(n46_adj_246), 
         .Z(n19)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut.init = 16'hfefc;
    LUT4 i5_4_lut_adj_376 (.A(\read_value[12]_adj_199 ), .B(n10_adj_334), 
         .C(n8_adj_200), .D(n32141), .Z(n13_adj_180)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_376.init = 16'hfefc;
    LUT4 Select_4285_i8_2_lut (.A(databus_out[1]), .B(rw), .Z(n8_adj_330)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4285_i8_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_377 (.A(\read_value[1]_adj_201 ), .B(n14_adj_337), 
         .C(n3_adj_202), .D(n32161), .Z(n18_adj_331)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_377.init = 16'hfefc;
    LUT4 i1_4_lut_adj_378 (.A(read_value_adj_288[1]), .B(read_value_adj_289[1]), 
         .C(n52_adj_129), .D(n64), .Z(n12_adj_332)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_378.init = 16'heca0;
    LUT4 i5_4_lut_adj_379 (.A(\read_value[1]_adj_203 ), .B(read_value_adj_287[1]), 
         .C(n32141), .D(n46), .Z(n16)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i5_4_lut_adj_379.init = 16'heca0;
    LUT4 i3_4_lut_adj_380 (.A(read_value[1]), .B(read_value_adj_290[1]), 
         .C(n52), .D(n19559), .Z(n14_adj_337)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_380.init = 16'heca0;
    LUT4 Select_4260_i5_2_lut (.A(databus_out[14]), .B(rw), .Z(n5_adj_318)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4260_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_381 (.A(read_value[14]), .B(\read_value[14]_adj_204 ), 
         .C(n52), .D(n32164), .Z(n10_adj_319)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_381.init = 16'heca0;
    LUT4 i3_4_lut_adj_382 (.A(read_value_adj_287[12]), .B(read_value_adj_288[12]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_181)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_382.init = 16'heca0;
    LUT4 i7_4_lut_adj_383 (.A(n13_adj_349), .B(n11_adj_350), .C(n2_adj_205), 
         .D(n5_adj_352), .Z(databus[9])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_383.init = 16'hfffe;
    LUT4 i5_4_lut_adj_384 (.A(\read_value[9]_adj_206 ), .B(n10_adj_179), 
         .C(n8_adj_207), .D(n32141), .Z(n13_adj_349)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_384.init = 16'hfefc;
    LUT4 i7_4_lut_adj_385 (.A(n13_adj_355), .B(n11_adj_356), .C(n2_adj_208), 
         .D(n5_adj_221), .Z(databus[13])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_385.init = 16'hfffe;
    LUT4 i5_4_lut_adj_386 (.A(\read_value[13]_adj_209 ), .B(n10_adj_287), 
         .C(n8_adj_210), .D(n32141), .Z(n13_adj_355)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_386.init = 16'hfefc;
    LUT4 i3_4_lut_adj_387 (.A(read_value_adj_287[9]), .B(read_value_adj_288[9]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_350)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_387.init = 16'heca0;
    LUT4 i3_4_lut_adj_388 (.A(read_value_adj_287[13]), .B(read_value_adj_288[13]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_356)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_388.init = 16'heca0;
    LUT4 Select_4227_i5_2_lut (.A(databus_out[25]), .B(n34064), .Z(n5_c)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4227_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_389 (.A(read_value[25]), .B(\read_value[25]_adj_211 ), 
         .C(n52), .D(n32164), .Z(n10_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_389.init = 16'heca0;
    LUT4 i3_4_lut_adj_390 (.A(read_value_adj_287[21]), .B(read_value_adj_288[21]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_368)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_390.init = 16'heca0;
    LUT4 Select_4275_i5_2_lut (.A(databus_out[9]), .B(n34064), .Z(n5_adj_352)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4275_i5_2_lut.init = 16'h2222;
    LUT4 n1150_bdd_3_lut_23642 (.A(n1150), .B(\register_addr[0] ), .C(\register[1] [3]), 
         .Z(n31833)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1150_bdd_3_lut_23642.init = 16'he2e2;
    LUT4 n1150_bdd_3_lut_23603 (.A(\register[2] [3]), .B(\register[3] [3]), 
         .C(\register_addr[0] ), .Z(n31832)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1150_bdd_3_lut_23603.init = 16'hcaca;
    LUT4 Select_4218_i5_2_lut (.A(databus_out[28]), .B(n34064), .Z(n5_adj_176)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4218_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_391 (.A(read_value[28]), .B(\read_value[28]_adj_212 ), 
         .C(n52), .D(n32164), .Z(n10_adj_270)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_391.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_23486 (.A(\register[6] [4]), .B(\register_addr[0] ), 
         .Z(n31575)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23486.init = 16'h2222;
    L6MUX21 i23723 (.D0(n32105), .D1(n32102), .SD(\register_addr[2] ), 
            .Z(n32106));
    LUT4 Select_4239_i5_2_lut (.A(databus_out[21]), .B(rw), .Z(n5_adj_371)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4239_i5_2_lut.init = 16'h2222;
    PFUMX i23721 (.BLUT(n32104), .ALUT(n32103), .C0(\register_addr[1] ), 
          .Z(n32105));
    LUT4 register_addr_1__bdd_2_lut_23453 (.A(\register[6] [6]), .B(\register_addr[0] ), 
         .Z(n31521)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_23453.init = 16'h2222;
    LUT4 i7_4_lut_adj_392 (.A(n13_adj_372), .B(n11_adj_373), .C(n2_adj_213), 
         .D(n5_adj_375), .Z(databus[27])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_392.init = 16'hfffe;
    LUT4 register_addr_1__bdd_3_lut_23454 (.A(\register_addr[0] ), .B(\register[4] [6]), 
         .C(\register[5] [6]), .Z(n31522)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23454.init = 16'he4e4;
    PFUMX i23719 (.BLUT(n32101), .ALUT(n32100), .C0(\register_addr[1] ), 
          .Z(n32102));
    LUT4 i5_4_lut_adj_393 (.A(\read_value[27]_adj_214 ), .B(n10_adj_376), 
         .C(n8_adj_215), .D(n32141), .Z(n13_adj_372)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_393.init = 16'hfefc;
    LUT4 i3_4_lut_adj_394 (.A(read_value_adj_287[27]), .B(read_value_adj_288[27]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_373)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_394.init = 16'heca0;
    LUT4 i14_2_lut (.A(\select[7] ), .B(n34064), .Z(n46_adj_246)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(214[19:32])
    defparam i14_2_lut.init = 16'h8888;
    LUT4 n1165_bdd_3_lut_23898 (.A(n1165), .B(\register_addr[0] ), .C(\register[1] [6]), 
         .Z(n31525)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1165_bdd_3_lut_23898.init = 16'he2e2;
    LUT4 Select_4221_i5_2_lut (.A(databus_out[27]), .B(n34064), .Z(n5_adj_375)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4221_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_395 (.A(read_value[27]), .B(\read_value[27]_adj_216 ), 
         .C(n52), .D(n32164), .Z(n10_adj_376)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_395.init = 16'heca0;
    LUT4 i2_4_lut_adj_396 (.A(read_value[21]), .B(\read_value[21]_adj_217 ), 
         .C(n52), .D(n32164), .Z(n10_adj_192)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_396.init = 16'heca0;
    L6MUX21 i23670 (.D0(n31986), .D1(n31983), .SD(\register_addr[2] ), 
            .Z(n31987));
    PFUMX i23668 (.BLUT(n31985), .ALUT(n31984), .C0(\register_addr[1] ), 
          .Z(n31986));
    LUT4 i10_4_lut_adj_397 (.A(n15_adj_384), .B(n20_adj_385), .C(n2_adj_218), 
         .D(n7_adj_387), .Z(databus[6])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_397.init = 16'hfffe;
    LUT4 i4_4_lut_adj_398 (.A(\read_value[6]_adj_219 ), .B(\read_value[6]_adj_220 ), 
         .C(n32164), .D(n32161), .Z(n15_adj_384)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_398.init = 16'heca0;
    PFUMX i23665 (.BLUT(n31982), .ALUT(n31981), .C0(\register_addr[1] ), 
          .Z(n31983));
    PFUMX i23413 (.BLUT(n31522), .ALUT(n31521), .C0(\register_addr[1] ), 
          .Z(n31523));
    L6MUX21 i23661 (.D0(n31979), .D1(n31976), .SD(\register_addr[2] ), 
            .Z(n31980));
    PFUMX i23656 (.BLUT(n31975), .ALUT(n31974), .C0(\register_addr[1] ), 
          .Z(n31976));
    LUT4 i7_4_lut_adj_399 (.A(n13_adj_389), .B(n11_adj_390), .C(n2_adj_221), 
         .D(n5_adj_392), .Z(databus[24])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_399.init = 16'hfffe;
    FD1S3IX read_value__i1 (.D(n31712), .CK(\select[7] ), .CD(n32185), 
            .Q(read_value_adj_556[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1S3IX read_value__i2 (.D(n31987), .CK(\select[7] ), .CD(n32185), 
            .Q(read_value_adj_556[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1S3IX read_value__i3 (.D(n31835), .CK(\select[7] ), .CD(n32185), 
            .Q(read_value_adj_556[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1S3IX read_value__i4 (.D(n31581), .CK(\select[7] ), .CD(n32185), 
            .Q(read_value_adj_556[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1S3IX read_value__i5 (.D(n32106), .CK(\select[7] ), .CD(n32185), 
            .Q(read_value_adj_556[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1S3IX read_value__i6 (.D(n31527), .CK(\select[7] ), .CD(n32185), 
            .Q(read_value_adj_556[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1S3IX read_value__i7 (.D(n31980), .CK(\select[7] ), .CD(n32185), 
            .Q(read_value_adj_556[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i7.GSR = "ENABLED";
    LUT4 i9_4_lut_adj_400 (.A(read_value_adj_556[6]), .B(n18_adj_395), .C(n12_adj_396), 
         .D(n46_adj_246), .Z(n20_adj_385)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_400.init = 16'hfefc;
    LUT4 register_addr_1__bdd_3_lut_23487 (.A(\register_addr[0] ), .B(\register[4] [4]), 
         .C(\register[5] [4]), .Z(n31576)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_23487.init = 16'he4e4;
    PFUMX i23659 (.BLUT(n31978), .ALUT(n31977), .C0(\register_addr[1] ), 
          .Z(n31979));
    LUT4 i5_4_lut_adj_401 (.A(\read_value[24]_adj_222 ), .B(n10_adj_397), 
         .C(n8_adj_223), .D(n32141), .Z(n13_adj_389)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_401.init = 16'hfefc;
    LUT4 i3_4_lut_adj_402 (.A(read_size[0]), .B(read_size_c[0]), .C(\select[1] ), 
         .D(\select[7] ), .Z(n13)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_402.init = 16'heca0;
    LUT4 i8_4_lut_adj_403 (.A(\read_size[0]_adj_224 ), .B(n16_adj_402), 
         .C(n9), .D(n32215), .Z(n18)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_403.init = 16'hfefc;
    LUT4 i4_4_lut_adj_404 (.A(\read_size[0]_adj_225 ), .B(\read_size[0]_adj_226 ), 
         .C(n32182), .D(\select[2] ), .Z(n14)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_404.init = 16'heca0;
    LUT4 i6_4_lut (.A(\read_size[0]_adj_227 ), .B(n12_adj_408), .C(n5), 
         .D(n32155), .Z(n16_adj_402)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut.init = 16'hfefc;
    LUT4 i2_4_lut_adj_405 (.A(\read_size[0]_adj_228 ), .B(\read_size[0]_adj_229 ), 
         .C(\select[5] ), .D(n32203), .Z(n12_adj_408)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_405.init = 16'heca0;
    LUT4 Select_4280_i7_2_lut (.A(databus_out[6]), .B(n34064), .Z(n7_adj_387)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4280_i7_2_lut.init = 16'h2222;
    LUT4 i3_4_lut_adj_406 (.A(n32178), .B(n6), .C(n1), .D(\read_size[2]_adj_230 ), 
         .Z(\reg_size[2] )) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_406.init = 16'hfefc;
    LUT4 i7_4_lut_adj_407 (.A(read_value_adj_287[6]), .B(n14_adj_414), .C(n3_adj_231), 
         .D(n46), .Z(n18_adj_395)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_407.init = 16'hfefc;
    LUT4 i2_4_lut_adj_408 (.A(\read_size[2]_adj_232 ), .B(n32), .C(n32182), 
         .D(n32251), .Z(n6)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_408.init = 16'heca0;
    LUT4 Select_4290_i1_2_lut (.A(read_size[2]), .B(\select[1] ), .Z(n1)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4290_i1_2_lut.init = 16'h8888;
    LUT4 i7_4_lut_adj_409 (.A(n13_adj_418), .B(n11_adj_419), .C(n2_adj_233), 
         .D(n5_adj_421), .Z(databus[26])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_409.init = 16'hfffe;
    LUT4 i5_4_lut_adj_410 (.A(\read_value[26]_adj_234 ), .B(n10_adj_422), 
         .C(n8_adj_235), .D(n32141), .Z(n13_adj_418)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_410.init = 16'hfefc;
    LUT4 i3_4_lut_adj_411 (.A(read_value_adj_287[24]), .B(read_value_adj_288[24]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_390)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_411.init = 16'heca0;
    LUT4 i3_4_lut_adj_412 (.A(read_value_adj_287[26]), .B(read_value_adj_288[26]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_419)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_412.init = 16'heca0;
    LUT4 Select_4224_i5_2_lut (.A(databus_out[26]), .B(n34064), .Z(n5_adj_421)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4224_i5_2_lut.init = 16'h2222;
    LUT4 Select_4230_i5_2_lut (.A(databus_out[24]), .B(rw), .Z(n5_adj_392)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4230_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_413 (.A(read_value[26]), .B(\read_value[26]_adj_236 ), 
         .C(n52), .D(n32164), .Z(n10_adj_422)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_413.init = 16'heca0;
    L6MUX21 i23630 (.D0(n31910), .D1(n31907), .SD(\register_addr[2] ), 
            .Z(n31911));
    PFUMX i23628 (.BLUT(n31909), .ALUT(n31908), .C0(\register_addr[1] ), 
          .Z(n31910));
    LUT4 i1_4_lut_adj_414 (.A(read_value_adj_288[6]), .B(read_value_adj_289[6]), 
         .C(n52_adj_129), .D(n64), .Z(n12_adj_396)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_414.init = 16'heca0;
    LUT4 i2_4_lut_adj_415 (.A(read_value[24]), .B(\read_value[24]_adj_237 ), 
         .C(n52), .D(n32164), .Z(n10_adj_397)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_415.init = 16'heca0;
    LUT4 i2_4_lut_adj_416 (.A(read_value[12]), .B(\read_value[12]_adj_238 ), 
         .C(n52), .D(n32164), .Z(n10_adj_334)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_416.init = 16'heca0;
    PFUMX i23625 (.BLUT(n31906), .ALUT(n31905), .C0(\register_addr[1] ), 
          .Z(n31907));
    LUT4 i10_4_lut_adj_417 (.A(n15_adj_436), .B(n20_adj_437), .C(n2_adj_239), 
         .D(n7_adj_439), .Z(databus[0])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_417.init = 16'hfffe;
    LUT4 i4_4_lut_adj_418 (.A(\read_value[0]_adj_240 ), .B(\read_value[0]_adj_241 ), 
         .C(n32164), .D(n32161), .Z(n15_adj_436)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_418.init = 16'heca0;
    LUT4 i9_4_lut_adj_419 (.A(read_value_adj_556[0]), .B(n18_adj_442), .C(n12_adj_443), 
         .D(n46_adj_246), .Z(n20_adj_437)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_419.init = 16'hfefc;
    FD1S3IX read_value__i0 (.D(n31911), .CK(\select[7] ), .CD(n32185), 
            .Q(read_value_adj_556[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=708, LSE_RLINE=720 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(217[9] 229[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 Select_4286_i7_2_lut (.A(databus_out[0]), .B(rw), .Z(n7_adj_439)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4286_i7_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_420 (.A(read_value_adj_287[0]), .B(n14_adj_445), .C(n3_adj_242), 
         .D(n46), .Z(n18_adj_442)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_420.init = 16'hfefc;
    L6MUX21 i23606 (.D0(n31834), .D1(n31831), .SD(\register_addr[2] ), 
            .Z(n31835));
    LUT4 i1_4_lut_adj_421 (.A(read_value_adj_288[0]), .B(read_value_adj_289[0]), 
         .C(n52_adj_129), .D(n64), .Z(n12_adj_443)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_421.init = 16'heca0;
    LUT4 i3_4_lut_adj_422 (.A(read_value[0]), .B(read_value_adj_290[0]), 
         .C(n52), .D(n19559), .Z(n14_adj_445)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_422.init = 16'heca0;
    PFUMX i23604 (.BLUT(n31833), .ALUT(n31832), .C0(\register_addr[1] ), 
          .Z(n31834));
    LUT4 i7_4_lut_adj_423 (.A(n13_adj_451), .B(n11_adj_452), .C(n2_adj_243), 
         .D(n5_adj_454), .Z(databus[31])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_423.init = 16'hfffe;
    LUT4 i5_4_lut_adj_424 (.A(\read_value[31]_adj_244 ), .B(n10_adj_455), 
         .C(n8_adj_245), .D(n32141), .Z(n13_adj_451)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_424.init = 16'hfefc;
    LUT4 i3_4_lut_adj_425 (.A(read_value_adj_287[31]), .B(read_value_adj_288[31]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_452)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_425.init = 16'heca0;
    LUT4 Select_4209_i5_2_lut (.A(databus_out[31]), .B(n34064), .Z(n5_adj_454)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4209_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_426 (.A(read_value[31]), .B(\read_value[31]_adj_246 ), 
         .C(n52), .D(n32164), .Z(n10_adj_455)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_426.init = 16'heca0;
    PFUMX i23601 (.BLUT(n31830), .ALUT(n31829), .C0(\register_addr[1] ), 
          .Z(n31831));
    LUT4 i10_4_lut_adj_427 (.A(n15_adj_461), .B(n20_adj_462), .C(n2_adj_247), 
         .D(n7_adj_464), .Z(databus[7])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_427.init = 16'hfffe;
    LUT4 i7_4_lut_adj_428 (.A(n13_adj_465), .B(n11_adj_466), .C(n2_adj_248), 
         .D(n5_adj_468), .Z(databus[23])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_428.init = 16'hfffe;
    LUT4 i10_4_lut_adj_429 (.A(n15_adj_469), .B(n20_adj_470), .C(n2_adj_249), 
         .D(n7), .Z(databus[4])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_429.init = 16'hfffe;
    LUT4 i3_4_lut_adj_430 (.A(read_value[6]), .B(n19559), .C(n52), .D(read_value_adj_290[6]), 
         .Z(n14_adj_414)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_430.init = 16'heca0;
    LUT4 i1_2_lut (.A(\register_addr[0] ), .B(\register_addr[1] ), .Z(n29920)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i7_4_lut_adj_431 (.A(n13_adj_474), .B(n11_adj_475), .C(n2_adj_250), 
         .D(n5_adj_477), .Z(databus[30])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_431.init = 16'hfffe;
    LUT4 i5_4_lut_adj_432 (.A(\read_value[30]_adj_251 ), .B(n10_adj_478), 
         .C(n8_adj_252), .D(n32141), .Z(n13_adj_474)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_432.init = 16'hfefc;
    LUT4 i3_4_lut_adj_433 (.A(read_value_adj_287[30]), .B(read_value_adj_288[30]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_475)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_433.init = 16'heca0;
    LUT4 Select_4212_i5_2_lut (.A(databus_out[30]), .B(rw), .Z(n5_adj_477)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4212_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_434 (.A(read_value[30]), .B(\read_value[30]_adj_253 ), 
         .C(n52), .D(n32164), .Z(n10_adj_478)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_434.init = 16'heca0;
    LUT4 i4_4_lut_adj_435 (.A(\read_value[7]_adj_254 ), .B(\read_value[7]_adj_255 ), 
         .C(n32164), .D(n32161), .Z(n15_adj_461)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_435.init = 16'heca0;
    LUT4 i7_4_lut_adj_436 (.A(n13_adj_486), .B(n11_adj_487), .C(n2_adj_256), 
         .D(n5_adj_489), .Z(databus[29])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_436.init = 16'hfffe;
    LUT4 i5_4_lut_adj_437 (.A(\read_value[29]_adj_257 ), .B(n10_adj_490), 
         .C(n8_adj_258), .D(n32141), .Z(n13_adj_486)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_437.init = 16'hfefc;
    LUT4 i3_4_lut_adj_438 (.A(read_value_adj_287[29]), .B(read_value_adj_288[29]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_487)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_438.init = 16'heca0;
    LUT4 Select_4215_i5_2_lut (.A(databus_out[29]), .B(rw), .Z(n5_adj_489)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4215_i5_2_lut.init = 16'h2222;
    L6MUX21 i23540 (.D0(n31711), .D1(n31708), .SD(\register_addr[2] ), 
            .Z(n31712));
    PFUMX i23538 (.BLUT(n31710), .ALUT(n31709), .C0(\register_addr[1] ), 
          .Z(n31711));
    LUT4 i2_4_lut_adj_439 (.A(read_value[29]), .B(\read_value[29]_adj_259 ), 
         .C(n52), .D(n32164), .Z(n10_adj_490)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_439.init = 16'heca0;
    LUT4 i9_4_lut_adj_440 (.A(read_value_adj_556[7]), .B(n18_adj_496), .C(n12_adj_497), 
         .D(n46_adj_246), .Z(n20_adj_462)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_440.init = 16'hfefc;
    LUT4 i4_4_lut_adj_441 (.A(\read_value[4]_adj_260 ), .B(\read_value[4]_adj_261 ), 
         .C(n32164), .D(n32161), .Z(n15_adj_469)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_441.init = 16'heca0;
    PFUMX i23535 (.BLUT(n31707), .ALUT(n31706), .C0(\register_addr[1] ), 
          .Z(n31708));
    LUT4 i10_4_lut_adj_442 (.A(n15_adj_500), .B(n20_adj_501), .C(n2_adj_262), 
         .D(n7_adj_503), .Z(databus[5])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut_adj_442.init = 16'hfffe;
    LUT4 i4_4_lut_adj_443 (.A(\read_value[5]_adj_263 ), .B(\read_value[5]_adj_264 ), 
         .C(n32164), .D(n32161), .Z(n15_adj_500)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_443.init = 16'heca0;
    LUT4 i9_4_lut_adj_444 (.A(read_value_adj_556[5]), .B(n18_adj_506), .C(n12_adj_507), 
         .D(n46_adj_246), .Z(n20_adj_501)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_444.init = 16'hfefc;
    LUT4 i5_4_lut_adj_445 (.A(\read_value[23]_adj_265 ), .B(n10_adj_508), 
         .C(n8_adj_266), .D(n32141), .Z(n13_adj_465)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_445.init = 16'hfefc;
    LUT4 i3_4_lut_adj_446 (.A(read_value_adj_287[23]), .B(read_value_adj_288[23]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_466)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_446.init = 16'heca0;
    LUT4 i9_4_lut_adj_447 (.A(read_value_adj_556[4]), .B(n18_c), .C(n12), 
         .D(n46_adj_246), .Z(n20_adj_470)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i9_4_lut_adj_447.init = 16'hfefc;
    LUT4 Select_4279_i7_2_lut (.A(databus_out[7]), .B(rw), .Z(n7_adj_464)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4279_i7_2_lut.init = 16'h2222;
    LUT4 Select_4281_i7_2_lut (.A(databus_out[5]), .B(n34064), .Z(n7_adj_503)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4281_i7_2_lut.init = 16'h2222;
    LUT4 Select_4233_i5_2_lut (.A(databus_out[23]), .B(n34064), .Z(n5_adj_468)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4233_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_448 (.A(read_value[23]), .B(\read_value[23]_adj_267 ), 
         .C(n52), .D(n32164), .Z(n10_adj_508)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_448.init = 16'heca0;
    LUT4 i7_4_lut_adj_449 (.A(read_value_adj_287[7]), .B(n14_adj_515), .C(n3_adj_268), 
         .D(n46), .Z(n18_adj_496)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_449.init = 16'hfefc;
    LUT4 i7_4_lut_adj_450 (.A(read_value_adj_287[5]), .B(n14_adj_518), .C(n3_adj_269), 
         .D(n46), .Z(n18_adj_506)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i7_4_lut_adj_450.init = 16'hfefc;
    LUT4 i7_4_lut_adj_451 (.A(n13_adj_520), .B(n11_adj_521), .C(n2_adj_270), 
         .D(n5_adj_523), .Z(databus[22])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_451.init = 16'hfffe;
    LUT4 i1_4_lut_adj_452 (.A(read_value_adj_288[7]), .B(read_value_adj_289[7]), 
         .C(n52_adj_129), .D(n64), .Z(n12_adj_497)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_452.init = 16'heca0;
    LUT4 i3_4_lut_adj_453 (.A(read_value[7]), .B(n19559), .C(n52), .D(read_value_adj_290[7]), 
         .Z(n14_adj_515)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_453.init = 16'heca0;
    LUT4 i5_4_lut_adj_454 (.A(\read_value[22]_adj_271 ), .B(n10_adj_528), 
         .C(n8_adj_272), .D(n32141), .Z(n13_adj_520)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_454.init = 16'hfefc;
    LUT4 i1_4_lut_adj_455 (.A(read_value_adj_288[5]), .B(read_value_adj_289[5]), 
         .C(n52_adj_129), .D(n64), .Z(n12_adj_507)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_455.init = 16'heca0;
    LUT4 i3_4_lut_adj_456 (.A(read_value[5]), .B(n19559), .C(n52), .D(read_value_adj_290[5]), 
         .Z(n14_adj_518)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_456.init = 16'heca0;
    LUT4 i3_4_lut_adj_457 (.A(read_value_adj_287[22]), .B(read_value_adj_288[22]), 
         .C(n46), .D(n52_adj_129), .Z(n11_adj_521)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_457.init = 16'heca0;
    LUT4 Select_4236_i5_2_lut (.A(databus_out[22]), .B(n34064), .Z(n5_adj_523)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_4236_i5_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_458 (.A(read_value[22]), .B(\read_value[22]_adj_273 ), 
         .C(n52), .D(n32164), .Z(n10_adj_528)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_458.init = 16'heca0;
    L6MUX21 i23459 (.D0(n31580), .D1(n31577), .SD(\register_addr[2] ), 
            .Z(n31581));
    PFUMX i23457 (.BLUT(n31579), .ALUT(n31578), .C0(\register_addr[1] ), 
          .Z(n31580));
    LUT4 i7_4_lut_adj_459 (.A(n13_adj_194), .B(n11_adj_368), .C(n2_adj_274), 
         .D(n5_adj_371), .Z(databus[21])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_459.init = 16'hfffe;
    PWMReceiver recv_ch8 (.\count[6] (\count[6] ), .\count[5] (\count[5] ), 
            .n29947(n29947), .n5(n5_adj_275), .GND_net(GND_net), .n30260(n30260), 
            .\count[8] (\count[8] ), .\count[9] (\count[9] ), .n30482(n30482), 
            .n32135(n32135), .n30304(n30304), .n32302(n32302), .\count[4] (\count[4] ), 
            .n32245(n32245), .n32301(n32301), .n28333(n28333), .debug_c_c(debug_c_c), 
            .rc_ch8_c(rc_ch8_c), .n32256(n32256), .\count[1] (\count[1] ), 
            .\count[2] (\count[2] ), .n32257(n32257), .\count[3] (\count[3] ), 
            .n32218(n32218), .n32258(n32258), .\register[6] ({\register[6] }), 
            .n13605(n13605), .\count[0] (\count[0] ), .n30001(n30001), 
            .n29948(n29948), .n28141(n28141), .n1180(n1180), .n28234(n28234), 
            .n32129(n32129)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(257[14] 261[36])
    PWMReceiver_U1 recv_ch7 (.GND_net(GND_net), .debug_c_c(debug_c_c), .n32135(n32135), 
            .\register[5] ({\register[5] }), .n32134(n32134), .n30474(n30474), 
            .rc_ch7_c(rc_ch7_c), .n30623(n30623), .n1165(n1165), .n28140(n28140)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(252[14] 256[36])
    PWMReceiver_U2 recv_ch4 (.n32283(n32283), .n28331(n28331), .n32317(n32317), 
            .debug_c_c(debug_c_c), .n32135(n32135), .GND_net(GND_net), 
            .\register[4] ({\register[4] }), .n13974(n13974), .rc_ch4_c(rc_ch4_c), 
            .n28133(n28133), .n30472(n30472), .n1150(n1150), .n28233(n28233)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(247[14] 251[36])
    PWMReceiver_U3 recv_ch3 (.n32221(n32221), .\count[9] (\count[9]_adj_276 ), 
            .n32264(n32264), .n28330(n28330), .n5(n5_adj_277), .\count[5] (\count[5]_adj_278 ), 
            .n5_adj_57(n5_adj_279), .\count[6] (\count[6]_adj_280 ), .n32267(n32267), 
            .debug_c_c(debug_c_c), .n32135(n32135), .GND_net(GND_net), 
            .\count[8] (\count[8]_adj_281 ), .\register[3] ({\register[3] }), 
            .n13975(n13975), .rc_ch3_c(rc_ch3_c), .n28132(n28132), .n1135(n1135), 
            .n28222(n28222), .n32127(n32127), .n30470(n30470), .n30302(n30302)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(242[14] 246[36])
    PWMReceiver_U4 recv_ch2 (.n1120(n1120), .debug_c_c(debug_c_c), .n28232(n28232), 
            .n32125(n32125), .n32294(n32294), .GND_net(GND_net), .\count[9] (\count[9]_adj_282 ), 
            .\count[8] (\count[8]_adj_283 ), .\count[5] (\count[5]_adj_284 ), 
            .\count[6] (\count[6]_adj_285 ), .n32135(n32135), .rc_ch2_c(rc_ch2_c), 
            .\register[2] ({\register[2] }), .n13976(n13976), .n5(n5_adj_286), 
            .n32293(n32293), .n41(n41), .n28329(n28329), .n32296(n32296), 
            .n28144(n28144), .n30308(n30308), .n30465(n30465)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(237[14] 241[36])
    PWMReceiver_U5 recv_ch1 (.\register[1] ({\register[1] }), .debug_c_c(debug_c_c), 
            .n13977(n13977), .n30463(n30463), .n32135(n32135), .GND_net(GND_net), 
            .n32274(n32274), .n28328(n28328), .n32308(n32308), .rc_ch1_c(rc_ch1_c), 
            .n1105(n1105), .n28231(n28231), .n28129(n28129)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(232[17] 236[36])
    
endmodule
//
// Verilog Description of module PWMReceiver
//

module PWMReceiver (\count[6] , \count[5] , n29947, n5, GND_net, n30260, 
            \count[8] , \count[9] , n30482, n32135, n30304, n32302, 
            \count[4] , n32245, n32301, n28333, debug_c_c, rc_ch8_c, 
            n32256, \count[1] , \count[2] , n32257, \count[3] , n32218, 
            n32258, \register[6] , n13605, \count[0] , n30001, n29948, 
            n28141, n1180, n28234, n32129) /* synthesis syn_module_defined=1 */ ;
    output \count[6] ;
    output \count[5] ;
    output n29947;
    output n5;
    input GND_net;
    output n30260;
    output \count[8] ;
    output \count[9] ;
    output n30482;
    input n32135;
    output n30304;
    input n32302;
    output \count[4] ;
    input n32245;
    output n32301;
    output n28333;
    input debug_c_c;
    input rc_ch8_c;
    output n32256;
    output \count[1] ;
    output \count[2] ;
    output n32257;
    output \count[3] ;
    output n32218;
    output n32258;
    output [7:0]\register[6] ;
    input n13605;
    output \count[0] ;
    input n30001;
    input n29948;
    output n28141;
    output n1180;
    input n28234;
    input n32129;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n1174, n1186, n27074;
    wire [15:0]n116;
    
    wire n27073, n27072, n32210, n22747, n27071, n54, n30089, 
        n4, n10, n24, n4_adj_171, n16753, n9;
    wire [7:0]n230;
    wire [7:0]n43;
    
    wire n32209, n32244, n32299, n12910, n13409, n32243, n28289, 
        n28055, n4_adj_172, n27070, n28273, n27069, n27068, n27067, 
        n27566, n27565, n27564, n27563, n30233, n29673;
    
    LUT4 i1_2_lut_3_lut (.A(count[7]), .B(\count[6] ), .C(\count[5] ), 
         .Z(n29947)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i5_2_lut (.A(n1174), .B(n1186), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    CCU2D add_1783_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27074), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_17.INIT0 = 16'hd222;
    defparam add_1783_17.INIT1 = 16'h0000;
    defparam add_1783_17.INJECT1_0 = "NO";
    defparam add_1783_17.INJECT1_1 = "NO";
    CCU2D add_1783_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27073), 
          .COUT(n27074), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_15.INIT0 = 16'hd222;
    defparam add_1783_15.INIT1 = 16'hd222;
    defparam add_1783_15.INJECT1_0 = "NO";
    defparam add_1783_15.INJECT1_1 = "NO";
    CCU2D add_1783_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27072), 
          .COUT(n27073), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_13.INIT0 = 16'hd222;
    defparam add_1783_13.INIT1 = 16'hd222;
    defparam add_1783_13.INJECT1_0 = "NO";
    defparam add_1783_13.INJECT1_1 = "NO";
    LUT4 i3_3_lut_rep_389 (.A(n30260), .B(\count[6] ), .C(\count[8] ), 
         .Z(n32210)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i3_3_lut_rep_389.init = 16'hfefe;
    LUT4 i16051_2_lut_4_lut (.A(n30260), .B(\count[6] ), .C(\count[8] ), 
         .D(\count[9] ), .Z(n22747)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i16051_2_lut_4_lut.init = 16'hfe00;
    CCU2D add_1783_11 (.A0(\count[9] ), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27071), 
          .COUT(n27072), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_11.INIT0 = 16'hd222;
    defparam add_1783_11.INIT1 = 16'hd222;
    defparam add_1783_11.INJECT1_0 = "NO";
    defparam add_1783_11.INJECT1_1 = "NO";
    LUT4 i23080_4_lut (.A(n54), .B(n30089), .C(n4), .D(n10), .Z(n30482)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i23080_4_lut.init = 16'h3323;
    LUT4 i2_4_lut (.A(n32135), .B(n30304), .C(n24), .D(n4_adj_171), 
         .Z(n16753)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut.init = 16'h2000;
    LUT4 i31_3_lut (.A(n9), .B(n32210), .C(\count[9] ), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i31_3_lut.init = 16'h3a3a;
    LUT4 i1_2_lut (.A(n1174), .B(n1186), .Z(n4_adj_171)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i15634_2_lut (.A(n230[7]), .B(n4), .Z(n43[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15634_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_311 (.A(n32209), .B(\count[8] ), .C(n32302), .D(n32244), 
         .Z(n4)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i2_4_lut_adj_311.init = 16'hfbbb;
    LUT4 i3_4_lut (.A(\count[4] ), .B(n32245), .C(\count[8] ), .D(n29947), 
         .Z(n9)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i22801_4_lut (.A(count[12]), .B(n32301), .C(count[13]), .D(n32299), 
         .Z(n30304)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22801_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_478 (.A(count[11]), .B(count[10]), .Z(n32299)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_478.init = 16'heeee;
    LUT4 i21_4_lut (.A(n12910), .B(n13409), .C(n22747), .D(n32299), 
         .Z(n54)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_rep_422_3_lut (.A(count[11]), .B(count[10]), .C(\count[9] ), 
         .Z(n32243)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_422_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_adj_312 (.A(n1186), .B(n1174), .Z(n30089)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_312.init = 16'hbbbb;
    LUT4 i15633_2_lut (.A(n230[6]), .B(n4), .Z(n43[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15633_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_rep_388_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(n13409), 
         .D(\count[9] ), .Z(n32209)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_388_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_480 (.A(count[15]), .B(count[14]), .Z(n32301)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_480.init = 16'heeee;
    LUT4 i2_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(count[12]), 
         .D(count[13]), .Z(n13409)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_4_lut_adj_313 (.A(count[15]), .B(count[14]), .C(n5), 
         .D(n28333), .Z(n28289)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_313.init = 16'hfffe;
    LUT4 i15632_2_lut (.A(n230[5]), .B(n4), .Z(n43[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15632_2_lut.init = 16'h2222;
    LUT4 i15631_2_lut (.A(n230[4]), .B(n4), .Z(n43[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15631_2_lut.init = 16'h2222;
    LUT4 i15630_2_lut (.A(n230[3]), .B(n4), .Z(n43[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15630_2_lut.init = 16'h2222;
    FD1P3AX prev_in_46 (.D(n1186), .SP(n32135), .CK(debug_c_c), .Q(n1174));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch8_c), .SP(n32135), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1186));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(\count[9] ), .B(n32299), .C(n9), .D(n13409), 
         .Z(n12910)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i15085_2_lut_rep_435 (.A(\count[4] ), .B(\count[5] ), .Z(n32256)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15085_2_lut_rep_435.init = 16'h8888;
    LUT4 i22757_3_lut_4_lut (.A(\count[4] ), .B(\count[5] ), .C(n28055), 
         .D(count[7]), .Z(n30260)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i22757_3_lut_4_lut.init = 16'hff80;
    LUT4 i3292_2_lut_rep_436 (.A(\count[1] ), .B(\count[2] ), .Z(n32257)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3292_2_lut_rep_436.init = 16'h8888;
    LUT4 i2_3_lut_rep_397_4_lut (.A(\count[1] ), .B(\count[2] ), .C(\count[3] ), 
         .D(\count[4] ), .Z(n32218)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i2_3_lut_rep_397_4_lut.init = 16'hfff8;
    LUT4 i1_3_lut_4_lut (.A(\count[1] ), .B(\count[2] ), .C(\count[3] ), 
         .D(\count[4] ), .Z(n4_adj_172)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i1_2_lut_rep_437 (.A(count[7]), .B(\count[6] ), .Z(n32258)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_437.init = 16'h8888;
    LUT4 i1_2_lut_rep_423_3_lut_4_lut (.A(count[7]), .B(\count[6] ), .C(\count[5] ), 
         .D(\count[4] ), .Z(n32244)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_423_3_lut_4_lut.init = 16'h8000;
    CCU2D add_1783_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(\count[8] ), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27070), 
          .COUT(n27071), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_9.INIT0 = 16'hd222;
    defparam add_1783_9.INIT1 = 16'hd222;
    defparam add_1783_9.INJECT1_0 = "NO";
    defparam add_1783_9.INJECT1_1 = "NO";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    LUT4 i15629_2_lut (.A(n230[2]), .B(n4), .Z(n43[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15629_2_lut.init = 16'h2222;
    LUT4 i15628_2_lut (.A(n230[1]), .B(n4), .Z(n43[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15628_2_lut.init = 16'h2222;
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(\count[9] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(\count[8] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(\count[6] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(\count[5] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(\count[4] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(\count[3] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(\count[2] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(\count[1] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n13605), .PD(n16753), .CK(debug_c_c), 
            .Q(\register[6] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n13605), .PD(n16753), .CK(debug_c_c), 
            .Q(\register[6] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n13605), .PD(n16753), .CK(debug_c_c), 
            .Q(\register[6] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n13605), .PD(n16753), .CK(debug_c_c), 
            .Q(\register[6] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n13605), .PD(n16753), .CK(debug_c_c), 
            .Q(\register[6] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n13605), .PD(n16753), .CK(debug_c_c), 
            .Q(\register[6] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n13605), .PD(n16753), .CK(debug_c_c), 
            .Q(\register[6] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_314 (.A(count[13]), .B(count[12]), .C(n28273), .D(n32243), 
         .Z(n28333)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_314.init = 16'h8880;
    LUT4 i2_4_lut_adj_315 (.A(n32258), .B(\count[5] ), .C(\count[8] ), 
         .D(n4_adj_172), .Z(n28273)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_315.init = 16'ha080;
    CCU2D add_1783_7 (.A0(\count[5] ), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(\count[6] ), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27069), 
          .COUT(n27070), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_7.INIT0 = 16'hd222;
    defparam add_1783_7.INIT1 = 16'hd222;
    defparam add_1783_7.INJECT1_0 = "NO";
    defparam add_1783_7.INJECT1_1 = "NO";
    CCU2D add_1783_5 (.A0(\count[3] ), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(\count[4] ), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27068), 
          .COUT(n27069), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_5.INIT0 = 16'hd222;
    defparam add_1783_5.INIT1 = 16'hd222;
    defparam add_1783_5.INJECT1_0 = "NO";
    defparam add_1783_5.INJECT1_1 = "NO";
    CCU2D add_1783_3 (.A0(\count[1] ), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(\count[2] ), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27067), 
          .COUT(n27068), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_3.INIT0 = 16'hd222;
    defparam add_1783_3.INIT1 = 16'hd222;
    defparam add_1783_3.INJECT1_0 = "NO";
    defparam add_1783_3.INJECT1_1 = "NO";
    CCU2D add_1783_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n28289), .B1(n1186), .C1(\count[0] ), .D1(n1174), .COUT(n27067), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1783_1.INIT0 = 16'hF000;
    defparam add_1783_1.INIT1 = 16'ha565;
    defparam add_1783_1.INJECT1_0 = "NO";
    defparam add_1783_1.INJECT1_1 = "NO";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(\count[0] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    CCU2D sub_51_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27566), 
          .S0(n230[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_9.INIT1 = 16'h0000;
    defparam sub_51_add_2_9.INJECT1_0 = "NO";
    defparam sub_51_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_7 (.A0(\count[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count[6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27565), .COUT(n27566), .S0(n230[5]), .S1(n230[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_7.INJECT1_0 = "NO";
    defparam sub_51_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_5 (.A0(\count[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count[4] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27564), .COUT(n27565), .S0(n230[3]), .S1(n230[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_5.INJECT1_0 = "NO";
    defparam sub_51_add_2_5.INJECT1_1 = "NO";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n13605), .PD(n16753), .CK(debug_c_c), 
            .Q(\register[6] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D sub_51_add_2_3 (.A0(\count[1] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count[2] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27563), .COUT(n27564), .S0(n230[1]), .S1(n230[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_3.INJECT1_0 = "NO";
    defparam sub_51_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count[0] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27563), .S1(n230[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_1.INIT0 = 16'hF000;
    defparam sub_51_add_2_1.INIT1 = 16'h5555;
    defparam sub_51_add_2_1.INJECT1_0 = "NO";
    defparam sub_51_add_2_1.INJECT1_1 = "NO";
    LUT4 i10_3_lut_4_lut (.A(\count[8] ), .B(n32209), .C(n30001), .D(n29948), 
         .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i10_3_lut_4_lut.init = 16'h0100;
    LUT4 i22733_3_lut_4_lut (.A(\count[8] ), .B(n32209), .C(n29948), .D(n30001), 
         .Z(n30233)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i22733_3_lut_4_lut.init = 16'hfeee;
    LUT4 i15077_2_lut (.A(n230[0]), .B(n4), .Z(n43[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15077_2_lut.init = 16'h2222;
    LUT4 i1_4_lut (.A(n30233), .B(n30089), .C(n32299), .D(n29673), .Z(n28141)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hcecc;
    LUT4 i3_4_lut_adj_316 (.A(n54), .B(n22747), .C(n4), .D(n13409), 
         .Z(n29673)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut_adj_316.init = 16'h0010;
    LUT4 i3_4_lut_adj_317 (.A(\count[0] ), .B(\count[1] ), .C(\count[2] ), 
         .D(\count[3] ), .Z(n28055)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_317.init = 16'hfffe;
    FD1P3AX valid_48 (.D(n32129), .SP(n28234), .CK(debug_c_c), .Q(n1180));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMReceiver_U1
//

module PWMReceiver_U1 (GND_net, debug_c_c, n32135, \register[5] , n32134, 
            n30474, rc_ch7_c, n30623, n1165, n28140) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    input n32135;
    output [7:0]\register[5] ;
    input n32134;
    output n30474;
    input rc_ch7_c;
    output n30623;
    output n1165;
    input n28140;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27075;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n32288;
    wire [15:0]n116;
    
    wire n27076, n30010, n1171, n1159, n32286, n4, n13288, n32214, 
        n4_adj_168, n32192, n32287, n32190, n4_adj_169, n32179, 
        n16899;
    wire [7:0]n43;
    
    wire n54, n30039, n10, n30192, n32191, n5, n6, n28038, n6_adj_170, 
        n13323, n30048, n27883;
    wire [7:0]n230;
    
    wire n30011, n30049, n30184, n28035, n28586, n30194, n27562, 
        n27561, n27560, n27559, n27082, n27081, n27080, n27079, 
        n27078, n27077;
    
    CCU2D add_1779_3 (.A0(count[1]), .B0(n32288), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n32288), .C1(GND_net), .D1(GND_net), .CIN(n27075), 
          .COUT(n27076), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_3.INIT0 = 16'hd222;
    defparam add_1779_3.INIT1 = 16'hd222;
    defparam add_1779_3.INJECT1_0 = "NO";
    defparam add_1779_3.INJECT1_1 = "NO";
    CCU2D add_1779_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n30010), .B1(n1171), .C1(count[0]), .D1(n1159), .COUT(n27075), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_1.INIT0 = 16'hF000;
    defparam add_1779_1.INIT1 = 16'ha565;
    defparam add_1779_1.INJECT1_0 = "NO";
    defparam add_1779_1.INJECT1_1 = "NO";
    LUT4 i3248_2_lut_rep_465 (.A(count[1]), .B(count[2]), .Z(n32286)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3248_2_lut_rep_465.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[1]), .B(count[2]), .C(count[3]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_393 (.A(count[9]), .B(n13288), .Z(n32214)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_393.init = 16'heeee;
    LUT4 i1_3_lut_rep_371_4_lut (.A(count[9]), .B(n13288), .C(n4_adj_168), 
         .D(count[8]), .Z(n32192)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_3_lut_rep_371_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_466 (.A(count[6]), .B(count[7]), .Z(n32287)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_rep_466.init = 16'h8888;
    LUT4 i1_2_lut_rep_369_3_lut (.A(count[9]), .B(n13288), .C(count[8]), 
         .Z(n32190)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_369_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_adj_303 (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n4_adj_169)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i1_2_lut_3_lut_adj_303.init = 16'h8080;
    LUT4 i5_2_lut_rep_467 (.A(n1159), .B(n1171), .Z(n32288)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_467.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_304 (.A(n1159), .B(n1171), .C(n32179), .Z(n30010)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i1_2_lut_3_lut_adj_304.init = 16'hf4f4;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n32134), .PD(n16899), .CK(debug_c_c), 
            .Q(\register[5] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n32134), .PD(n16899), .CK(debug_c_c), 
            .Q(\register[5] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n32134), .PD(n16899), .CK(debug_c_c), 
            .Q(\register[5] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n32134), .PD(n16899), .CK(debug_c_c), 
            .Q(\register[5] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n32134), .PD(n16899), .CK(debug_c_c), 
            .Q(\register[5] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n32134), .PD(n16899), .CK(debug_c_c), 
            .Q(\register[5] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n32134), .PD(n16899), .CK(debug_c_c), 
            .Q(\register[5] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i23072_4_lut (.A(n54), .B(n30039), .C(n32192), .D(n10), .Z(n30474)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i23072_4_lut.init = 16'h3332;
    LUT4 i21_4_lut (.A(count[8]), .B(n30192), .C(n32214), .D(n32191), 
         .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h3230;
    LUT4 i22694_4_lut (.A(n13288), .B(count[9]), .C(n5), .D(n6), .Z(n30192)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i22694_4_lut.init = 16'heeea;
    LUT4 i2_2_lut (.A(count[7]), .B(count[8]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3_4_lut (.A(count[2]), .B(count[3]), .C(count[1]), .D(count[0]), 
         .Z(n28038)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut (.A(count[1]), .B(count[3]), .C(n6_adj_170), .D(n32287), 
         .Z(n4_adj_168)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'h8000;
    LUT4 i3_4_lut_adj_305 (.A(count[13]), .B(n13323), .C(count[12]), .D(n30048), 
         .Z(n13288)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_305.init = 16'hfffe;
    LUT4 i2_4_lut (.A(count[5]), .B(count[4]), .C(n32287), .D(n4), .Z(n27883)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut.init = 16'ha080;
    LUT4 i1_2_lut (.A(n1171), .B(n1159), .Z(n30039)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    FD1P3AX prev_in_46 (.D(n1171), .SP(n32135), .CK(debug_c_c), .Q(n1159));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch7_c), .SP(n32135), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1171));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut (.A(count[5]), .B(count[4]), .C(n28038), .D(count[6]), 
         .Z(n5)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i2_2_lut_3_lut (.A(count[5]), .B(count[4]), .C(count[2]), .Z(n6_adj_170)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_2_lut_3_lut.init = 16'h8080;
    LUT4 i15623_2_lut_4_lut (.A(count[8]), .B(n32214), .C(n4_adj_168), 
         .D(n230[3]), .Z(n43[3])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15623_2_lut_4_lut.init = 16'h0200;
    LUT4 i15622_2_lut_4_lut (.A(count[8]), .B(n32214), .C(n4_adj_168), 
         .D(n230[2]), .Z(n43[2])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15622_2_lut_4_lut.init = 16'h0200;
    LUT4 i10183_2_lut_3_lut (.A(n32135), .B(n30474), .C(n54), .Z(n16899)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i10183_2_lut_3_lut.init = 16'h8080;
    LUT4 i23234_3_lut_3_lut_4_lut (.A(n27883), .B(n32190), .C(n30192), 
         .D(n32179), .Z(n30011)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i23234_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i15621_2_lut_4_lut (.A(count[8]), .B(n32214), .C(n4_adj_168), 
         .D(n230[1]), .Z(n43[1])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15621_2_lut_4_lut.init = 16'h0200;
    LUT4 i1_4_lut_rep_358 (.A(n13323), .B(count[13]), .C(count[12]), .D(n30049), 
         .Z(n32179)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_rep_358.init = 16'heaaa;
    LUT4 i15074_2_lut_4_lut (.A(count[8]), .B(n32214), .C(n4_adj_168), 
         .D(n230[0]), .Z(n43[0])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15074_2_lut_4_lut.init = 16'h0200;
    LUT4 i22686_2_lut_4_lut (.A(count[8]), .B(n32214), .C(n4_adj_168), 
         .D(n54), .Z(n30184)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (D)) */ ;
    defparam i22686_2_lut_4_lut.init = 16'hff02;
    LUT4 i2_4_lut_adj_306 (.A(n30048), .B(count[9]), .C(n28035), .D(n4_adj_169), 
         .Z(n30049)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_306.init = 16'hfeee;
    LUT4 i2_4_lut_adj_307 (.A(count[5]), .B(count[4]), .C(n32286), .D(count[3]), 
         .Z(n28035)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    defparam i2_4_lut_adj_307.init = 16'hfeee;
    LUT4 i1_2_lut_adj_308 (.A(count[10]), .B(count[11]), .Z(n30048)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_308.init = 16'heeee;
    LUT4 i1_2_lut_adj_309 (.A(count[15]), .B(count[14]), .Z(n13323)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_309.init = 16'heeee;
    LUT4 i23221_4_lut (.A(n28586), .B(n32288), .C(n32179), .D(n30039), 
         .Z(n30623)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i23221_4_lut.init = 16'h3031;
    LUT4 i5_4_lut (.A(n30192), .B(n30184), .C(n32190), .D(n30194), .Z(n28586)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i5_4_lut.init = 16'h1110;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n32134), .PD(n16899), .CK(debug_c_c), 
            .Q(\register[5] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D sub_51_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27562), 
          .S0(n230[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_9.INIT1 = 16'h0000;
    defparam sub_51_add_2_9.INJECT1_0 = "NO";
    defparam sub_51_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27561), 
          .COUT(n27562), .S0(n230[5]), .S1(n230[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_7.INJECT1_0 = "NO";
    defparam sub_51_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27560), 
          .COUT(n27561), .S0(n230[3]), .S1(n230[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_5.INJECT1_0 = "NO";
    defparam sub_51_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27559), 
          .COUT(n27560), .S0(n230[1]), .S1(n230[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_3.INJECT1_0 = "NO";
    defparam sub_51_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27559), 
          .S1(n230[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_1.INIT0 = 16'hF000;
    defparam sub_51_add_2_1.INIT1 = 16'h5555;
    defparam sub_51_add_2_1.INJECT1_0 = "NO";
    defparam sub_51_add_2_1.INJECT1_1 = "NO";
    CCU2D add_1779_17 (.A0(count[15]), .B0(n32288), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27082), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_17.INIT0 = 16'hd222;
    defparam add_1779_17.INIT1 = 16'h0000;
    defparam add_1779_17.INJECT1_0 = "NO";
    defparam add_1779_17.INJECT1_1 = "NO";
    CCU2D add_1779_15 (.A0(count[13]), .B0(n32288), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n32288), .C1(GND_net), .D1(GND_net), .CIN(n27081), 
          .COUT(n27082), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_15.INIT0 = 16'hd222;
    defparam add_1779_15.INIT1 = 16'hd222;
    defparam add_1779_15.INJECT1_0 = "NO";
    defparam add_1779_15.INJECT1_1 = "NO";
    CCU2D add_1779_13 (.A0(count[11]), .B0(n32288), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n32288), .C1(GND_net), .D1(GND_net), .CIN(n27080), 
          .COUT(n27081), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_13.INIT0 = 16'hd222;
    defparam add_1779_13.INIT1 = 16'hd222;
    defparam add_1779_13.INJECT1_0 = "NO";
    defparam add_1779_13.INJECT1_1 = "NO";
    CCU2D add_1779_11 (.A0(count[9]), .B0(n32288), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n32288), .C1(GND_net), .D1(GND_net), .CIN(n27079), 
          .COUT(n27080), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_11.INIT0 = 16'hd222;
    defparam add_1779_11.INIT1 = 16'hd222;
    defparam add_1779_11.INJECT1_0 = "NO";
    defparam add_1779_11.INJECT1_1 = "NO";
    CCU2D add_1779_9 (.A0(count[7]), .B0(n32288), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n32288), .C1(GND_net), .D1(GND_net), .CIN(n27078), 
          .COUT(n27079), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_9.INIT0 = 16'hd222;
    defparam add_1779_9.INIT1 = 16'hd222;
    defparam add_1779_9.INJECT1_0 = "NO";
    defparam add_1779_9.INJECT1_1 = "NO";
    CCU2D add_1779_7 (.A0(count[5]), .B0(n32288), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n32288), .C1(GND_net), .D1(GND_net), .CIN(n27077), 
          .COUT(n27078), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_7.INIT0 = 16'hd222;
    defparam add_1779_7.INIT1 = 16'hd222;
    defparam add_1779_7.INJECT1_0 = "NO";
    defparam add_1779_7.INJECT1_1 = "NO";
    CCU2D add_1779_5 (.A0(count[3]), .B0(n32288), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n32288), .C1(GND_net), .D1(GND_net), .CIN(n27076), 
          .COUT(n27077), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1779_5.INIT0 = 16'hd222;
    defparam add_1779_5.INIT1 = 16'hd222;
    defparam add_1779_5.INJECT1_0 = "NO";
    defparam add_1779_5.INJECT1_1 = "NO";
    FD1P3AX valid_48 (.D(n30011), .SP(n28140), .CK(debug_c_c), .Q(n1165));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n32214), .C(n32191), 
         .D(n27883), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2_2_lut_rep_370 (.A(count[0]), .B(n4_adj_168), .Z(n32191)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_rep_370.init = 16'h8888;
    LUT4 i2_2_lut_3_lut_adj_310 (.A(count[0]), .B(n4_adj_168), .C(n27883), 
         .Z(n30194)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_310.init = 16'h8080;
    LUT4 i15627_2_lut_4_lut (.A(count[8]), .B(n32214), .C(n4_adj_168), 
         .D(n230[7]), .Z(n43[7])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15627_2_lut_4_lut.init = 16'h0200;
    LUT4 i15625_2_lut_4_lut (.A(count[8]), .B(n32214), .C(n4_adj_168), 
         .D(n230[5]), .Z(n43[5])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15625_2_lut_4_lut.init = 16'h0200;
    LUT4 i15624_2_lut_4_lut (.A(count[8]), .B(n32214), .C(n4_adj_168), 
         .D(n230[4]), .Z(n43[4])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15624_2_lut_4_lut.init = 16'h0200;
    LUT4 i15626_2_lut_4_lut (.A(count[8]), .B(n32214), .C(n4_adj_168), 
         .D(n230[6]), .Z(n43[6])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i15626_2_lut_4_lut.init = 16'h0200;
    
endmodule
//
// Verilog Description of module PWMReceiver_U2
//

module PWMReceiver_U2 (n32283, n28331, n32317, debug_c_c, n32135, 
            GND_net, \register[4] , n13974, rc_ch4_c, n28133, n30472, 
            n1150, n28233) /* synthesis syn_module_defined=1 */ ;
    output n32283;
    output n28331;
    output n32317;
    input debug_c_c;
    input n32135;
    input GND_net;
    output [7:0]\register[4] ;
    input n13974;
    input rc_ch4_c;
    output n28133;
    output n30472;
    output n1150;
    input n28233;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n32259, n28189, n5, n32255, n41, n32260, n29791, n27857, 
        n32254;
    wire [7:0]n230;
    
    wire n4;
    wire [7:0]n43;
    
    wire n9, n32318, n32193, n30162, n54, n28201, n1144, n1156, 
        n28285;
    wire [15:0]n116;
    
    wire n16504, n32217, n30068, n30286, n44_adj_167, n30322, n32126, 
        n30004, n10, n30235, n30220, n29671, n24, n27090, n27089, 
        n27088, n27087, n27086, n27085, n27084, n27083, n27558, 
        n27557, n27556, n27555, n29792;
    
    LUT4 i15299_2_lut_rep_438 (.A(count[4]), .B(count[5]), .Z(n32259)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15299_2_lut_rep_438.init = 16'h8888;
    LUT4 i1_3_lut_4_lut (.A(count[4]), .B(count[5]), .C(count[7]), .D(n28189), 
         .Z(n5)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i2965_2_lut_rep_434_3_lut (.A(count[1]), .B(count[2]), .C(count[3]), 
         .Z(n32255)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2965_2_lut_rep_434_3_lut.init = 16'h8080;
    LUT4 i1_3_lut_4_lut_adj_295 (.A(count[1]), .B(count[2]), .C(count[4]), 
         .D(count[3]), .Z(n41)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i1_3_lut_4_lut_adj_295.init = 16'hfff8;
    LUT4 i1_2_lut_rep_439 (.A(count[7]), .B(count[6]), .Z(n32260)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_439.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[7]), .B(count[6]), .C(count[8]), .Z(n29791)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i2_3_lut_4_lut (.A(count[7]), .B(count[6]), .C(n41), .D(count[5]), 
         .Z(n27857)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_433_3_lut_4_lut (.A(count[7]), .B(count[6]), .C(count[5]), 
         .D(count[4]), .Z(n32254)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_433_3_lut_4_lut.init = 16'h8000;
    LUT4 i15068_2_lut (.A(n230[0]), .B(n4), .Z(n43[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15068_2_lut.init = 16'h2222;
    LUT4 i21_4_lut (.A(n9), .B(n32318), .C(n32193), .D(n30162), .Z(n54)) /* synthesis lut_function=(!(A (B+(D))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h0032;
    LUT4 i3_3_lut (.A(n5), .B(count[6]), .C(count[8]), .Z(n28201)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i3_3_lut.init = 16'hfefe;
    LUT4 i15619_2_lut (.A(n230[6]), .B(n4), .Z(n43[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15619_2_lut.init = 16'h2222;
    LUT4 i15618_2_lut (.A(n230[5]), .B(n4), .Z(n43[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15618_2_lut.init = 16'h2222;
    LUT4 i15617_2_lut (.A(n230[4]), .B(n4), .Z(n43[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15617_2_lut.init = 16'h2222;
    LUT4 i5_2_lut_rep_462 (.A(n1144), .B(n1156), .Z(n32283)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_462.init = 16'h4444;
    LUT4 i2_3_lut_4_lut_adj_296 (.A(n1144), .B(n1156), .C(n28331), .D(n32317), 
         .Z(n28285)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i2_3_lut_4_lut_adj_296.init = 16'hfff4;
    LUT4 i15616_2_lut (.A(n230[3]), .B(n4), .Z(n43[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15616_2_lut.init = 16'h2222;
    LUT4 i15615_2_lut (.A(n230[2]), .B(n4), .Z(n43[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15615_2_lut.init = 16'h2222;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    LUT4 i15614_2_lut (.A(n230[1]), .B(n4), .Z(n43[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15614_2_lut.init = 16'h2222;
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n13974), .PD(n16504), .CK(debug_c_c), 
            .Q(\register[4] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n13974), .PD(n16504), .CK(debug_c_c), 
            .Q(\register[4] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n13974), .PD(n16504), .CK(debug_c_c), 
            .Q(\register[4] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n13974), .PD(n16504), .CK(debug_c_c), 
            .Q(\register[4] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n13974), .PD(n16504), .CK(debug_c_c), 
            .Q(\register[4] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n13974), .PD(n16504), .CK(debug_c_c), 
            .Q(\register[4] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n13974), .PD(n16504), .CK(debug_c_c), 
            .Q(\register[4] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i3_3_lut_4_lut (.A(count[0]), .B(n32255), .C(n29791), .D(n32259), 
         .Z(n9)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_3_lut_4_lut.init = 16'h8000;
    LUT4 i22666_3_lut_4_lut (.A(count[13]), .B(n32217), .C(count[9]), 
         .D(n28201), .Z(n30162)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i22666_3_lut_4_lut.init = 16'hfeee;
    LUT4 i1_2_lut_rep_372_3_lut_4_lut (.A(n32317), .B(count[12]), .C(n30068), 
         .D(count[13]), .Z(n32193)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_372_3_lut_4_lut.init = 16'hfffe;
    LUT4 i22783_3_lut_4_lut (.A(n32317), .B(count[12]), .C(n32318), .D(count[13]), 
         .Z(n30286)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22783_3_lut_4_lut.init = 16'hfffe;
    LUT4 n44_bdd_4_lut (.A(n44_adj_167), .B(n30322), .C(count[9]), .D(n30286), 
         .Z(n32126)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n44_bdd_4_lut.init = 16'h00ca;
    FD1P3AX prev_in_46 (.D(n1156), .SP(n32135), .CK(debug_c_c), .Q(n1144));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch4_c), .SP(n32135), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1156));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_496 (.A(count[15]), .B(count[14]), .Z(n32317)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_496.init = 16'heeee;
    LUT4 i22763_2_lut_rep_396_3_lut (.A(count[15]), .B(count[14]), .C(count[12]), 
         .Z(n32217)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22763_2_lut_rep_396_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_497 (.A(count[11]), .B(count[10]), .Z(n32318)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_497.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_297 (.A(count[11]), .B(count[10]), .C(count[9]), 
         .Z(n30068)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_3_lut_adj_297.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32259), .B(n32260), .C(n32255), .D(count[0]), 
         .Z(n30004)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i10_3_lut_4_lut (.A(count[8]), .B(n32193), .C(n30004), .D(n27857), 
         .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i10_3_lut_4_lut.init = 16'h0100;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    LUT4 i22734_3_lut_4_lut (.A(count[8]), .B(n32193), .C(n27857), .D(n30004), 
         .Z(n30235)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i22734_3_lut_4_lut.init = 16'hfeee;
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n13974), .PD(n16504), .CK(debug_c_c), 
            .Q(\register[4] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n30235), .B(n30220), .C(n32318), .D(n29671), .Z(n28133)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hcecc;
    LUT4 i23070_4_lut (.A(n54), .B(n30220), .C(n4), .D(n10), .Z(n30472)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i23070_4_lut.init = 16'h3323;
    LUT4 i2_4_lut (.A(n32135), .B(n30286), .C(n24), .D(n30220), .Z(n16504)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut.init = 16'h0020;
    LUT4 i3_3_lut_adj_298 (.A(n54), .B(n30162), .C(n4), .Z(n29671)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i3_3_lut_adj_298.init = 16'h1010;
    LUT4 i31_3_lut (.A(n9), .B(n28201), .C(count[9]), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i31_3_lut.init = 16'h3a3a;
    LUT4 i15620_2_lut (.A(n230[7]), .B(n4), .Z(n43[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15620_2_lut.init = 16'h2222;
    CCU2D add_1775_17 (.A0(count[15]), .B0(n32283), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27090), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_17.INIT0 = 16'hd222;
    defparam add_1775_17.INIT1 = 16'h0000;
    defparam add_1775_17.INJECT1_0 = "NO";
    defparam add_1775_17.INJECT1_1 = "NO";
    CCU2D add_1775_15 (.A0(count[13]), .B0(n32283), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n32283), .C1(GND_net), .D1(GND_net), .CIN(n27089), 
          .COUT(n27090), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_15.INIT0 = 16'hd222;
    defparam add_1775_15.INIT1 = 16'hd222;
    defparam add_1775_15.INJECT1_0 = "NO";
    defparam add_1775_15.INJECT1_1 = "NO";
    CCU2D add_1775_13 (.A0(count[11]), .B0(n32283), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n32283), .C1(GND_net), .D1(GND_net), .CIN(n27088), 
          .COUT(n27089), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_13.INIT0 = 16'hd222;
    defparam add_1775_13.INIT1 = 16'hd222;
    defparam add_1775_13.INJECT1_0 = "NO";
    defparam add_1775_13.INJECT1_1 = "NO";
    CCU2D add_1775_11 (.A0(count[9]), .B0(n32283), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n32283), .C1(GND_net), .D1(GND_net), .CIN(n27087), 
          .COUT(n27088), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_11.INIT0 = 16'hd222;
    defparam add_1775_11.INIT1 = 16'hd222;
    defparam add_1775_11.INJECT1_0 = "NO";
    defparam add_1775_11.INJECT1_1 = "NO";
    CCU2D add_1775_9 (.A0(count[7]), .B0(n32283), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n32283), .C1(GND_net), .D1(GND_net), .CIN(n27086), 
          .COUT(n27087), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_9.INIT0 = 16'hd222;
    defparam add_1775_9.INIT1 = 16'hd222;
    defparam add_1775_9.INJECT1_0 = "NO";
    defparam add_1775_9.INJECT1_1 = "NO";
    CCU2D add_1775_7 (.A0(count[5]), .B0(n32283), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n32283), .C1(GND_net), .D1(GND_net), .CIN(n27085), 
          .COUT(n27086), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_7.INIT0 = 16'hd222;
    defparam add_1775_7.INIT1 = 16'hd222;
    defparam add_1775_7.INJECT1_0 = "NO";
    defparam add_1775_7.INJECT1_1 = "NO";
    CCU2D add_1775_5 (.A0(count[3]), .B0(n32283), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n32283), .C1(GND_net), .D1(GND_net), .CIN(n27084), 
          .COUT(n27085), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_5.INIT0 = 16'hd222;
    defparam add_1775_5.INIT1 = 16'hd222;
    defparam add_1775_5.INJECT1_0 = "NO";
    defparam add_1775_5.INJECT1_1 = "NO";
    CCU2D add_1775_3 (.A0(count[1]), .B0(n32283), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n32283), .C1(GND_net), .D1(GND_net), .CIN(n27083), 
          .COUT(n27084), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_3.INIT0 = 16'hd222;
    defparam add_1775_3.INIT1 = 16'hd222;
    defparam add_1775_3.INJECT1_0 = "NO";
    defparam add_1775_3.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_299 (.A(n32193), .B(count[8]), .C(n32255), .D(n32254), 
         .Z(n4)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i2_4_lut_adj_299.init = 16'hfbbb;
    CCU2D sub_51_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27558), 
          .S0(n230[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_9.INIT1 = 16'h0000;
    defparam sub_51_add_2_9.INJECT1_0 = "NO";
    defparam sub_51_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27557), 
          .COUT(n27558), .S0(n230[5]), .S1(n230[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_7.INJECT1_0 = "NO";
    defparam sub_51_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27556), 
          .COUT(n27557), .S0(n230[3]), .S1(n230[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_5.INJECT1_0 = "NO";
    defparam sub_51_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27555), 
          .COUT(n27556), .S0(n230[1]), .S1(n230[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_3.INJECT1_0 = "NO";
    defparam sub_51_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27555), 
          .S1(n230[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_1.INIT0 = 16'hF000;
    defparam sub_51_add_2_1.INIT1 = 16'h5555;
    defparam sub_51_add_2_1.INJECT1_0 = "NO";
    defparam sub_51_add_2_1.INJECT1_1 = "NO";
    CCU2D add_1775_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n28285), .B1(n1156), .C1(count[0]), .D1(n1144), .COUT(n27083), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1775_1.INIT0 = 16'hF000;
    defparam add_1775_1.INIT1 = 16'ha565;
    defparam add_1775_1.INJECT1_0 = "NO";
    defparam add_1775_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_300 (.A(count[8]), .B(n32260), .C(count[5]), .D(n41), 
         .Z(n44_adj_167)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_adj_300.init = 16'heaaa;
    LUT4 i23157_3_lut (.A(count[8]), .B(count[6]), .C(n5), .Z(n30322)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i23157_3_lut.init = 16'h0101;
    LUT4 i22721_2_lut (.A(n1144), .B(n1156), .Z(n30220)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i22721_2_lut.init = 16'hdddd;
    LUT4 i3_4_lut (.A(count[0]), .B(count[1]), .C(count[2]), .D(count[3]), 
         .Z(n28189)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    FD1P3AX valid_48 (.D(n32126), .SP(n28233), .CK(debug_c_c), .Q(n1150));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_301 (.A(count[13]), .B(count[12]), .C(n29792), .D(n30068), 
         .Z(n28331)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_301.init = 16'h8880;
    LUT4 i1_4_lut_adj_302 (.A(count[5]), .B(n29791), .C(count[4]), .D(n32255), 
         .Z(n29792)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_302.init = 16'hccc8;
    
endmodule
//
// Verilog Description of module PWMReceiver_U3
//

module PWMReceiver_U3 (n32221, \count[9] , n32264, n28330, n5, \count[5] , 
            n5_adj_57, \count[6] , n32267, debug_c_c, n32135, GND_net, 
            \count[8] , \register[3] , n13975, rc_ch3_c, n28132, n1135, 
            n28222, n32127, n30470, n30302) /* synthesis syn_module_defined=1 */ ;
    output n32221;
    output \count[9] ;
    output n32264;
    output n28330;
    output n5;
    output \count[5] ;
    output n5_adj_57;
    output \count[6] ;
    output n32267;
    input debug_c_c;
    input n32135;
    input GND_net;
    output \count[8] ;
    output [7:0]\register[3] ;
    input n13975;
    input rc_ch3_c;
    output n28132;
    output n1135;
    input n28222;
    input n32127;
    output n30470;
    output n30302;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n12959, n13403, n22701, n32263, n54;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n32262, n4;
    wire [7:0]n230;
    
    wire n4_adj_165;
    wire [7:0]n43;
    
    wire n32220, n32195, n28286, n32265, n32222, n32266, n28054, 
        n29899, n32219;
    wire [15:0]n116;
    
    wire n16507, n9, n29900, n29916, n1129, n1141, n30237, n30036, 
        n29669, n32196, n27098, n27097, n27096, n27095, n27094, 
        n27093, n27092, n27091, n28275, n10, n27554, n27553, n27552, 
        n27551, n24;
    
    LUT4 i21_4_lut (.A(n12959), .B(n13403), .C(n22701), .D(n32263), 
         .Z(n54)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h0002;
    LUT4 i3160_2_lut_rep_441 (.A(count[1]), .B(count[2]), .Z(n32262)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3160_2_lut_rep_441.init = 16'h8888;
    LUT4 i2_3_lut_rep_400_4_lut (.A(count[1]), .B(count[2]), .C(count[3]), 
         .D(count[4]), .Z(n32221)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i2_3_lut_rep_400_4_lut.init = 16'hfff8;
    LUT4 i1_3_lut_4_lut (.A(count[1]), .B(count[2]), .C(count[3]), .D(count[4]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i15063_2_lut (.A(n230[0]), .B(n4_adj_165), .Z(n43[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15063_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_rep_442 (.A(count[11]), .B(count[10]), .Z(n32263)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_442.init = 16'heeee;
    LUT4 i1_2_lut_rep_399_3_lut (.A(count[11]), .B(count[10]), .C(\count[9] ), 
         .Z(n32220)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_399_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_374_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(n13403), 
         .D(\count[9] ), .Z(n32195)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_374_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_443 (.A(count[15]), .B(count[14]), .Z(n32264)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_443.init = 16'heeee;
    LUT4 i2_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(count[12]), 
         .D(count[13]), .Z(n13403)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_4_lut_adj_287 (.A(count[15]), .B(count[14]), .C(n28330), 
         .D(n5), .Z(n28286)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_287.init = 16'hfffe;
    LUT4 i2_3_lut_rep_444 (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n32265)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_rep_444.init = 16'h8080;
    LUT4 i1_2_lut_rep_401_4_lut (.A(count[2]), .B(count[3]), .C(count[1]), 
         .D(count[0]), .Z(n32222)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_401_4_lut.init = 16'h8000;
    LUT4 i15477_2_lut_rep_445 (.A(count[4]), .B(\count[5] ), .Z(n32266)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15477_2_lut_rep_445.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_288 (.A(count[4]), .B(\count[5] ), .C(count[7]), 
         .D(n28054), .Z(n5_adj_57)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut_adj_288.init = 16'hf8f0;
    LUT4 i1_2_lut_rep_446 (.A(count[7]), .B(\count[6] ), .Z(n32267)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_446.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[7]), .B(\count[6] ), .C(\count[5] ), 
         .Z(n29899)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_398_3_lut_4_lut (.A(count[7]), .B(\count[6] ), .C(\count[5] ), 
         .D(count[4]), .Z(n32219)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_398_3_lut_4_lut.init = 16'h8000;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(\count[9] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(\count[8] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(\count[6] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(\count[5] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n13975), .PD(n16507), .CK(debug_c_c), 
            .Q(\register[3] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n13975), .PD(n16507), .CK(debug_c_c), 
            .Q(\register[3] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n13975), .PD(n16507), .CK(debug_c_c), 
            .Q(\register[3] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n13975), .PD(n16507), .CK(debug_c_c), 
            .Q(\register[3] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n13975), .PD(n16507), .CK(debug_c_c), 
            .Q(\register[3] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n13975), .PD(n16507), .CK(debug_c_c), 
            .Q(\register[3] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n13975), .PD(n16507), .CK(debug_c_c), 
            .Q(\register[3] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(\count[9] ), .B(n32263), .C(n9), .D(n13403), 
         .Z(n12959)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut (.A(count[4]), .B(count[3]), .C(n32262), .D(n29899), 
         .Z(n29900)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfe00;
    LUT4 i1_2_lut_3_lut_4_lut_adj_289 (.A(count[0]), .B(n32265), .C(n32267), 
         .D(n32266), .Z(n29916)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_289.init = 16'h8000;
    FD1P3AX prev_in_46 (.D(n1141), .SP(n32135), .CK(debug_c_c), .Q(n1129));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch3_c), .SP(n32135), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1141));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(n32195), .B(\count[8] ), .C(n32219), .D(n32265), 
         .Z(n4_adj_165)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i2_4_lut.init = 16'hfbbb;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n13975), .PD(n16507), .CK(debug_c_c), 
            .Q(\register[3] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i15612_2_lut (.A(n230[6]), .B(n4_adj_165), .Z(n43[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15612_2_lut.init = 16'h2222;
    LUT4 i1_4_lut (.A(n30237), .B(n30036), .C(n32263), .D(n29669), .Z(n28132)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hcecc;
    LUT4 i3_4_lut (.A(n54), .B(n13403), .C(n4_adj_165), .D(n22701), 
         .Z(n29669)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut.init = 16'h0010;
    LUT4 i3_3_lut_rep_375 (.A(n5_adj_57), .B(\count[6] ), .C(\count[8] ), 
         .Z(n32196)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i3_3_lut_rep_375.init = 16'hfefe;
    LUT4 i16005_2_lut_4_lut (.A(n5_adj_57), .B(\count[6] ), .C(\count[8] ), 
         .D(\count[9] ), .Z(n22701)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i16005_2_lut_4_lut.init = 16'hfe00;
    LUT4 i15611_2_lut (.A(n230[5]), .B(n4_adj_165), .Z(n43[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15611_2_lut.init = 16'h2222;
    LUT4 i15610_2_lut (.A(n230[4]), .B(n4_adj_165), .Z(n43[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15610_2_lut.init = 16'h2222;
    LUT4 i15609_2_lut (.A(n230[3]), .B(n4_adj_165), .Z(n43[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15609_2_lut.init = 16'h2222;
    LUT4 i5_2_lut (.A(n1129), .B(n1141), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut.init = 16'h4444;
    CCU2D add_1771_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27098), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1771_17.INIT0 = 16'hd222;
    defparam add_1771_17.INIT1 = 16'h0000;
    defparam add_1771_17.INJECT1_0 = "NO";
    defparam add_1771_17.INJECT1_1 = "NO";
    CCU2D add_1771_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27097), 
          .COUT(n27098), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1771_15.INIT0 = 16'hd222;
    defparam add_1771_15.INIT1 = 16'hd222;
    defparam add_1771_15.INJECT1_0 = "NO";
    defparam add_1771_15.INJECT1_1 = "NO";
    CCU2D add_1771_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27096), 
          .COUT(n27097), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1771_13.INIT0 = 16'hd222;
    defparam add_1771_13.INIT1 = 16'hd222;
    defparam add_1771_13.INJECT1_0 = "NO";
    defparam add_1771_13.INJECT1_1 = "NO";
    CCU2D add_1771_11 (.A0(\count[9] ), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27095), 
          .COUT(n27096), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1771_11.INIT0 = 16'hd222;
    defparam add_1771_11.INIT1 = 16'hd222;
    defparam add_1771_11.INJECT1_0 = "NO";
    defparam add_1771_11.INJECT1_1 = "NO";
    CCU2D add_1771_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(\count[8] ), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27094), 
          .COUT(n27095), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1771_9.INIT0 = 16'hd222;
    defparam add_1771_9.INIT1 = 16'hd222;
    defparam add_1771_9.INJECT1_0 = "NO";
    defparam add_1771_9.INJECT1_1 = "NO";
    CCU2D add_1771_7 (.A0(\count[5] ), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(\count[6] ), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27093), 
          .COUT(n27094), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1771_7.INIT0 = 16'hd222;
    defparam add_1771_7.INIT1 = 16'hd222;
    defparam add_1771_7.INJECT1_0 = "NO";
    defparam add_1771_7.INJECT1_1 = "NO";
    CCU2D add_1771_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27092), 
          .COUT(n27093), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1771_5.INIT0 = 16'hd222;
    defparam add_1771_5.INIT1 = 16'hd222;
    defparam add_1771_5.INJECT1_0 = "NO";
    defparam add_1771_5.INJECT1_1 = "NO";
    CCU2D add_1771_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27091), 
          .COUT(n27092), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1771_3.INIT0 = 16'hd222;
    defparam add_1771_3.INIT1 = 16'hd222;
    defparam add_1771_3.INJECT1_0 = "NO";
    defparam add_1771_3.INJECT1_1 = "NO";
    CCU2D add_1771_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n28286), .B1(n1141), .C1(count[0]), .D1(n1129), .COUT(n27091), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1771_1.INIT0 = 16'hF000;
    defparam add_1771_1.INIT1 = 16'ha565;
    defparam add_1771_1.INJECT1_0 = "NO";
    defparam add_1771_1.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_290 (.A(count[13]), .B(count[12]), .C(n28275), .D(n32220), 
         .Z(n28330)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_290.init = 16'h8880;
    LUT4 i2_4_lut_adj_291 (.A(n32267), .B(\count[5] ), .C(\count[8] ), 
         .D(n4), .Z(n28275)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_291.init = 16'ha080;
    LUT4 i10_3_lut_4_lut (.A(\count[8] ), .B(n32195), .C(n29916), .D(n29900), 
         .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i10_3_lut_4_lut.init = 16'h0100;
    LUT4 i22735_3_lut_4_lut (.A(\count[8] ), .B(n32195), .C(n29900), .D(n29916), 
         .Z(n30237)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i22735_3_lut_4_lut.init = 16'hfeee;
    LUT4 i15608_2_lut (.A(n230[2]), .B(n4_adj_165), .Z(n43[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15608_2_lut.init = 16'h2222;
    CCU2D sub_51_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27554), 
          .S0(n230[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_9.INIT1 = 16'h0000;
    defparam sub_51_add_2_9.INJECT1_0 = "NO";
    defparam sub_51_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_7 (.A0(\count[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count[6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27553), .COUT(n27554), .S0(n230[5]), .S1(n230[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_7.INJECT1_0 = "NO";
    defparam sub_51_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27552), 
          .COUT(n27553), .S0(n230[3]), .S1(n230[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_5.INJECT1_0 = "NO";
    defparam sub_51_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27551), 
          .COUT(n27552), .S0(n230[1]), .S1(n230[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_3.INJECT1_0 = "NO";
    defparam sub_51_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27551), 
          .S1(n230[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_1.INIT0 = 16'hF000;
    defparam sub_51_add_2_1.INIT1 = 16'h5555;
    defparam sub_51_add_2_1.INJECT1_0 = "NO";
    defparam sub_51_add_2_1.INJECT1_1 = "NO";
    FD1P3AX valid_48 (.D(n32127), .SP(n28222), .CK(debug_c_c), .Q(n1135));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i23068_4_lut (.A(n54), .B(n30036), .C(n4_adj_165), .D(n10), 
         .Z(n30470)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i23068_4_lut.init = 16'h3323;
    LUT4 i2_4_lut_adj_292 (.A(n32135), .B(n30302), .C(n24), .D(n30036), 
         .Z(n16507)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut_adj_292.init = 16'h0020;
    LUT4 i15607_2_lut (.A(n230[1]), .B(n4_adj_165), .Z(n43[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15607_2_lut.init = 16'h2222;
    LUT4 i31_3_lut (.A(n9), .B(n32196), .C(\count[9] ), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i31_3_lut.init = 16'h3a3a;
    LUT4 i15613_2_lut (.A(n230[7]), .B(n4_adj_165), .Z(n43[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15613_2_lut.init = 16'h2222;
    LUT4 i22799_4_lut (.A(count[12]), .B(n32264), .C(count[13]), .D(n32263), 
         .Z(n30302)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22799_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(n1141), .B(n1129), .Z(n30036)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i3_4_lut_adj_293 (.A(count[4]), .B(n32222), .C(\count[8] ), .D(n29899), 
         .Z(n9)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut_adj_293.init = 16'h8000;
    LUT4 i3_4_lut_adj_294 (.A(count[0]), .B(count[1]), .C(count[2]), .D(count[3]), 
         .Z(n28054)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_294.init = 16'hfffe;
    
endmodule
//
// Verilog Description of module PWMReceiver_U4
//

module PWMReceiver_U4 (n1120, debug_c_c, n28232, n32125, n32294, GND_net, 
            \count[9] , \count[8] , \count[5] , \count[6] , n32135, 
            rc_ch2_c, \register[2] , n13976, n5, n32293, n41, n28329, 
            n32296, n28144, n30308, n30465) /* synthesis syn_module_defined=1 */ ;
    output n1120;
    input debug_c_c;
    input n28232;
    input n32125;
    output n32294;
    input GND_net;
    output \count[9] ;
    output \count[8] ;
    output \count[5] ;
    output \count[6] ;
    input n32135;
    input rc_ch2_c;
    output [7:0]\register[2] ;
    input n13976;
    output n5;
    output n32293;
    output n41;
    output n28329;
    output n32296;
    output n28144;
    output n30308;
    output n30465;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27106;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    wire [15:0]n116;
    wire [7:0]n230;
    
    wire n4;
    wire [7:0]n43;
    
    wire n27105, n27104, n27103, n27102, n27101, n1126, n16509, 
        n32206, n32184, n32238, n29789, n30006, n30182, n27100, 
        n32240, n1114, n28359, n28200, n32295, n13397, n32207, 
        n32237, n32297, n32208, n4_adj_163, n30030, n12, n8, n32183, 
        n54, n9, n4_adj_164, n32186, n28274, n27099, n10, n24, 
        n27550, n27549, n27548, n27547;
    
    FD1P3AX valid_48 (.D(n32125), .SP(n28232), .CK(debug_c_c), .Q(n1120));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    CCU2D add_1767_17 (.A0(count[15]), .B0(n32294), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27106), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1767_17.INIT0 = 16'hd222;
    defparam add_1767_17.INIT1 = 16'h0000;
    defparam add_1767_17.INJECT1_0 = "NO";
    defparam add_1767_17.INJECT1_1 = "NO";
    LUT4 i15060_2_lut (.A(n230[0]), .B(n4), .Z(n43[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15060_2_lut.init = 16'h2222;
    CCU2D add_1767_15 (.A0(count[13]), .B0(n32294), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n32294), .C1(GND_net), .D1(GND_net), .CIN(n27105), 
          .COUT(n27106), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1767_15.INIT0 = 16'hd222;
    defparam add_1767_15.INIT1 = 16'hd222;
    defparam add_1767_15.INJECT1_0 = "NO";
    defparam add_1767_15.INJECT1_1 = "NO";
    CCU2D add_1767_13 (.A0(count[11]), .B0(n32294), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n32294), .C1(GND_net), .D1(GND_net), .CIN(n27104), 
          .COUT(n27105), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1767_13.INIT0 = 16'hd222;
    defparam add_1767_13.INIT1 = 16'hd222;
    defparam add_1767_13.INJECT1_0 = "NO";
    defparam add_1767_13.INJECT1_1 = "NO";
    CCU2D add_1767_11 (.A0(\count[9] ), .B0(n32294), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n32294), .C1(GND_net), .D1(GND_net), .CIN(n27103), 
          .COUT(n27104), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1767_11.INIT0 = 16'hd222;
    defparam add_1767_11.INIT1 = 16'hd222;
    defparam add_1767_11.INJECT1_0 = "NO";
    defparam add_1767_11.INJECT1_1 = "NO";
    CCU2D add_1767_9 (.A0(count[7]), .B0(n32294), .C0(GND_net), .D0(GND_net), 
          .A1(\count[8] ), .B1(n32294), .C1(GND_net), .D1(GND_net), 
          .CIN(n27102), .COUT(n27103), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1767_9.INIT0 = 16'hd222;
    defparam add_1767_9.INIT1 = 16'hd222;
    defparam add_1767_9.INJECT1_0 = "NO";
    defparam add_1767_9.INJECT1_1 = "NO";
    CCU2D add_1767_7 (.A0(\count[5] ), .B0(n32294), .C0(GND_net), .D0(GND_net), 
          .A1(\count[6] ), .B1(n32294), .C1(GND_net), .D1(GND_net), 
          .CIN(n27101), .COUT(n27102), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1767_7.INIT0 = 16'hd222;
    defparam add_1767_7.INIT1 = 16'hd222;
    defparam add_1767_7.INJECT1_0 = "NO";
    defparam add_1767_7.INJECT1_1 = "NO";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch2_c), .SP(n32135), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1126));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(\count[9] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(\count[8] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(\count[6] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(\count[5] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n13976), .PD(n16509), .CK(debug_c_c), 
            .Q(\register[2] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n13976), .PD(n16509), .CK(debug_c_c), 
            .Q(\register[2] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n13976), .PD(n16509), .CK(debug_c_c), 
            .Q(\register[2] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n13976), .PD(n16509), .CK(debug_c_c), 
            .Q(\register[2] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n13976), .PD(n16509), .CK(debug_c_c), 
            .Q(\register[2] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n13976), .PD(n16509), .CK(debug_c_c), 
            .Q(\register[2] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n13976), .PD(n16509), .CK(debug_c_c), 
            .Q(\register[2] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i3_3_lut_rep_385 (.A(n5), .B(\count[6] ), .C(\count[8] ), .Z(n32206)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i3_3_lut_rep_385.init = 16'hfefe;
    LUT4 i15852_2_lut_rep_363_4_lut (.A(n5), .B(\count[6] ), .C(\count[8] ), 
         .D(\count[9] ), .Z(n32184)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i15852_2_lut_rep_363_4_lut.init = 16'hfe00;
    LUT4 i2_2_lut_3_lut_4_lut (.A(count[0]), .B(n32238), .C(n29789), .D(n30006), 
         .Z(n30182)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_2_lut_3_lut_4_lut.init = 16'h8000;
    CCU2D add_1767_5 (.A0(count[3]), .B0(n32294), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n32294), .C1(GND_net), .D1(GND_net), .CIN(n27100), 
          .COUT(n27101), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1767_5.INIT0 = 16'hd222;
    defparam add_1767_5.INIT1 = 16'hd222;
    defparam add_1767_5.INJECT1_0 = "NO";
    defparam add_1767_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_472 (.A(count[7]), .B(\count[6] ), .Z(n32293)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_472.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[7]), .B(\count[6] ), .C(n41), 
         .D(\count[5] ), .Z(n29789)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_419_3_lut (.A(count[7]), .B(\count[6] ), .C(\count[5] ), 
         .Z(n32240)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_419_3_lut.init = 16'h8080;
    LUT4 i5_2_lut_rep_473 (.A(n1114), .B(n1126), .Z(n32294)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_473.init = 16'h4444;
    LUT4 i2_3_lut_4_lut (.A(n1114), .B(n1126), .C(n28329), .D(n32296), 
         .Z(n28359)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i2_3_lut_4_lut.init = 16'hfff4;
    LUT4 i1_3_lut_4_lut (.A(count[4]), .B(\count[5] ), .C(count[7]), .D(n28200), 
         .Z(n5)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_278 (.A(count[4]), .B(\count[5] ), .C(\count[6] ), 
         .D(count[7]), .Z(n30006)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_278.init = 16'h8000;
    LUT4 i1_2_lut_rep_474 (.A(count[11]), .B(count[10]), .Z(n32295)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_474.init = 16'heeee;
    LUT4 i1_2_lut_rep_386_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(n13397), 
         .D(\count[9] ), .Z(n32207)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_386_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_416_3_lut (.A(count[11]), .B(count[10]), .C(\count[9] ), 
         .Z(n32237)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_rep_416_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_475 (.A(count[15]), .B(count[14]), .Z(n32296)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_475.init = 16'heeee;
    LUT4 i2_3_lut_4_lut_adj_279 (.A(count[15]), .B(count[14]), .C(count[12]), 
         .D(count[13]), .Z(n13397)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_279.init = 16'hfffe;
    LUT4 i3116_2_lut_rep_476 (.A(count[1]), .B(count[2]), .Z(n32297)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3116_2_lut_rep_476.init = 16'h8888;
    LUT4 i2905_2_lut_rep_417_3_lut (.A(count[1]), .B(count[2]), .C(count[3]), 
         .Z(n32238)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2905_2_lut_rep_417_3_lut.init = 16'h8080;
    LUT4 i1_3_lut_4_lut_adj_280 (.A(count[1]), .B(count[2]), .C(count[4]), 
         .D(count[3]), .Z(n41)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i1_3_lut_4_lut_adj_280.init = 16'hfff8;
    LUT4 i1_2_lut_rep_387_3_lut_4_lut (.A(count[1]), .B(count[2]), .C(count[0]), 
         .D(count[3]), .Z(n32208)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_387_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_281 (.A(count[1]), .B(count[2]), .C(count[4]), 
         .D(count[3]), .Z(n4_adj_163)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_281.init = 16'hf8f0;
    LUT4 i1_4_lut (.A(n32184), .B(n30030), .C(n12), .D(n8), .Z(n28144)) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hdccc;
    LUT4 i5_4_lut (.A(n32183), .B(n13397), .C(n30182), .D(n32295), .Z(n12)) /* synthesis lut_function=(!(A (B+(D))+!A (B+((D)+!C)))) */ ;
    defparam i5_4_lut.init = 16'h0032;
    LUT4 i1_2_lut (.A(n54), .B(n4), .Z(n8)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i22805_4_lut (.A(count[12]), .B(n32296), .C(count[13]), .D(n32295), 
         .Z(n30308)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22805_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(n9), .B(n32295), .C(n32207), .D(n4_adj_164), 
         .Z(n54)) /* synthesis lut_function=(!(A (B+(D))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h0032;
    LUT4 i2_4_lut (.A(n32207), .B(\count[8] ), .C(n32238), .D(n30006), 
         .Z(n4)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i2_4_lut.init = 16'hfbbb;
    LUT4 i3_4_lut (.A(count[4]), .B(n32208), .C(\count[8] ), .D(n32240), 
         .Z(n9)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_362_3_lut_4_lut (.A(\count[9] ), .B(n32295), .C(\count[8] ), 
         .D(n13397), .Z(n32183)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_362_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_365_3_lut_4_lut (.A(n32297), .B(count[3]), .C(n30006), 
         .D(count[0]), .Z(n32186)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_365_3_lut_4_lut.init = 16'h8000;
    LUT4 i3_4_lut_adj_282 (.A(count[0]), .B(count[1]), .C(count[2]), .D(count[3]), 
         .Z(n28200)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_282.init = 16'hfffe;
    LUT4 i1_2_lut_adj_283 (.A(n1126), .B(n1114), .Z(n30030)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_283.init = 16'hbbbb;
    LUT4 i2_4_lut_adj_284 (.A(count[13]), .B(count[12]), .C(n28274), .D(n32237), 
         .Z(n28329)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_284.init = 16'h8880;
    LUT4 i2_4_lut_adj_285 (.A(n32293), .B(\count[5] ), .C(\count[8] ), 
         .D(n4_adj_163), .Z(n28274)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_285.init = 16'ha080;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n13976), .PD(n16509), .CK(debug_c_c), 
            .Q(\register[2] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D add_1767_3 (.A0(count[1]), .B0(n32294), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n32294), .C1(GND_net), .D1(GND_net), .CIN(n27099), 
          .COUT(n27100), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1767_3.INIT0 = 16'hd222;
    defparam add_1767_3.INIT1 = 16'hd222;
    defparam add_1767_3.INJECT1_0 = "NO";
    defparam add_1767_3.INJECT1_1 = "NO";
    FD1P3AX prev_in_46 (.D(n1126), .SP(n32135), .CK(debug_c_c), .Q(n1114));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    CCU2D add_1767_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n28359), .B1(n1126), .C1(count[0]), .D1(n1114), .COUT(n27099), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1767_1.INIT0 = 16'hF000;
    defparam add_1767_1.INIT1 = 16'ha565;
    defparam add_1767_1.INJECT1_0 = "NO";
    defparam add_1767_1.INJECT1_1 = "NO";
    LUT4 i23063_4_lut (.A(n54), .B(n30030), .C(n4), .D(n10), .Z(n30465)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i23063_4_lut.init = 16'h3323;
    LUT4 i2_4_lut_adj_286 (.A(n32135), .B(n30308), .C(n24), .D(n30030), 
         .Z(n16509)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut_adj_286.init = 16'h0020;
    LUT4 i31_3_lut (.A(n9), .B(n32206), .C(\count[9] ), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i31_3_lut.init = 16'h3a3a;
    LUT4 i15604_2_lut (.A(n230[7]), .B(n4), .Z(n43[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15604_2_lut.init = 16'h2222;
    LUT4 i10_3_lut_4_lut (.A(\count[8] ), .B(n32207), .C(n32186), .D(n29789), 
         .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i10_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_3_lut (.A(n32206), .B(\count[9] ), .C(n13397), .Z(n4_adj_164)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i15603_2_lut (.A(n230[6]), .B(n4), .Z(n43[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15603_2_lut.init = 16'h2222;
    LUT4 i15602_2_lut (.A(n230[5]), .B(n4), .Z(n43[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15602_2_lut.init = 16'h2222;
    LUT4 i15601_2_lut (.A(n230[4]), .B(n4), .Z(n43[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15601_2_lut.init = 16'h2222;
    LUT4 i15600_2_lut (.A(n230[3]), .B(n4), .Z(n43[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15600_2_lut.init = 16'h2222;
    LUT4 i15599_2_lut (.A(n230[2]), .B(n4), .Z(n43[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15599_2_lut.init = 16'h2222;
    LUT4 i15598_2_lut (.A(n230[1]), .B(n4), .Z(n43[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15598_2_lut.init = 16'h2222;
    CCU2D sub_51_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27550), 
          .S0(n230[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_9.INIT1 = 16'h0000;
    defparam sub_51_add_2_9.INJECT1_0 = "NO";
    defparam sub_51_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_7 (.A0(\count[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count[6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27549), .COUT(n27550), .S0(n230[5]), .S1(n230[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_7.INJECT1_0 = "NO";
    defparam sub_51_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27548), 
          .COUT(n27549), .S0(n230[3]), .S1(n230[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_5.INJECT1_0 = "NO";
    defparam sub_51_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27547), 
          .COUT(n27548), .S0(n230[1]), .S1(n230[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_3.INJECT1_0 = "NO";
    defparam sub_51_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27547), 
          .S1(n230[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_1.INIT0 = 16'hF000;
    defparam sub_51_add_2_1.INIT1 = 16'h5555;
    defparam sub_51_add_2_1.INJECT1_0 = "NO";
    defparam sub_51_add_2_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U5
//

module PWMReceiver_U5 (\register[1] , debug_c_c, n13977, n30463, n32135, 
            GND_net, n32274, n28328, n32308, rc_ch1_c, n1105, n28231, 
            n28129) /* synthesis syn_module_defined=1 */ ;
    output [7:0]\register[1] ;
    input debug_c_c;
    input n13977;
    output n30463;
    input n32135;
    input GND_net;
    output n32274;
    output n28328;
    output n32308;
    input rc_ch1_c;
    output n1105;
    input n28231;
    output n28129;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [7:0]n230;
    
    wire n4;
    wire [7:0]n43;
    
    wire n16511, n54, n30033, n10, n30334, n24, n9, n32212;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(133[16:21])
    
    wire n32188, n32248, n32312, n32250, n29785, n28191;
    wire [15:0]n116;
    
    wire n1099, n1111, n28288, n12914, n32211, n22550, n32309, 
        n32249, n32246, n5, n44_adj_161, n30318, n32124, n32307, 
        n32247, n4_adj_162, n32311, n32313, n29913, n29786, n30239, 
        n27546, n27545, n27544, n27543, n27114, n27113, n27112, 
        n27111, n27110, n27109, n27108, n29667, n28276, n27107;
    
    LUT4 i15053_2_lut (.A(n230[0]), .B(n4), .Z(n43[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15053_2_lut.init = 16'h2222;
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n13977), .PD(n16511), .CK(debug_c_c), 
            .Q(\register[1] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n13977), .PD(n16511), .CK(debug_c_c), 
            .Q(\register[1] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n13977), .PD(n16511), .CK(debug_c_c), 
            .Q(\register[1] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n13977), .PD(n16511), .CK(debug_c_c), 
            .Q(\register[1] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n13977), .PD(n16511), .CK(debug_c_c), 
            .Q(\register[1] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n13977), .PD(n16511), .CK(debug_c_c), 
            .Q(\register[1] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n13977), .PD(n16511), .CK(debug_c_c), 
            .Q(\register[1] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i23061_4_lut (.A(n54), .B(n30033), .C(n4), .D(n10), .Z(n30463)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i23061_4_lut.init = 16'h3323;
    LUT4 i2_4_lut (.A(n32135), .B(n30334), .C(n24), .D(n30033), .Z(n16511)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i2_4_lut.init = 16'h0020;
    LUT4 i31_3_lut (.A(n9), .B(n32212), .C(count[9]), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i31_3_lut.init = 16'h3a3a;
    LUT4 i15597_2_lut (.A(n230[7]), .B(n4), .Z(n43[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15597_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_270 (.A(n32188), .B(count[8]), .C(n32248), .D(n32312), 
         .Z(n4)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i2_4_lut_adj_270.init = 16'hfbbb;
    LUT4 i3_4_lut (.A(count[4]), .B(n32250), .C(count[8]), .D(n29785), 
         .Z(n9)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i3_4_lut_adj_271 (.A(count[0]), .B(count[1]), .C(count[2]), .D(count[3]), 
         .Z(n28191)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_271.init = 16'hfffe;
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i4.GSR = "ENABLED";
    LUT4 i5_2_lut_rep_453 (.A(n1099), .B(n1111), .Z(n32274)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i5_2_lut_rep_453.init = 16'h4444;
    LUT4 i2_3_lut_4_lut (.A(n1099), .B(n1111), .C(n28328), .D(n32308), 
         .Z(n28288)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(152[10:31])
    defparam i2_3_lut_4_lut.init = 16'hfff4;
    LUT4 i1_2_lut (.A(n1111), .B(n1099), .Z(n30033)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i21_4_lut (.A(n12914), .B(n32211), .C(n22550), .D(n32309), 
         .Z(n54)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[13:39])
    defparam i21_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[13]), .B(n32249), .C(n9), .D(n32246), 
         .Z(n12914)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[28:39])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i3_3_lut_rep_391 (.A(n5), .B(count[6]), .C(count[8]), .Z(n32212)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i3_3_lut_rep_391.init = 16'hfefe;
    LUT4 i15858_2_lut_4_lut (.A(n5), .B(count[6]), .C(count[8]), .D(count[9]), 
         .Z(n22550)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i15858_2_lut_4_lut.init = 16'hfe00;
    LUT4 n44_bdd_4_lut (.A(n44_adj_161), .B(n30318), .C(count[9]), .D(n30334), 
         .Z(n32124)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n44_bdd_4_lut.init = 16'h00ca;
    LUT4 i15596_2_lut (.A(n230[6]), .B(n4), .Z(n43[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15596_2_lut.init = 16'h2222;
    LUT4 i15595_2_lut (.A(n230[5]), .B(n4), .Z(n43[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15595_2_lut.init = 16'h2222;
    LUT4 i15594_2_lut (.A(n230[4]), .B(n4), .Z(n43[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15594_2_lut.init = 16'h2222;
    LUT4 i3072_2_lut_rep_486 (.A(count[1]), .B(count[2]), .Z(n32307)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3072_2_lut_rep_486.init = 16'h8888;
    LUT4 i2_3_lut_rep_426_4_lut (.A(count[1]), .B(count[2]), .C(count[3]), 
         .D(count[4]), .Z(n32247)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i2_3_lut_rep_426_4_lut.init = 16'hfff8;
    LUT4 i1_3_lut_4_lut (.A(count[1]), .B(count[2]), .C(count[3]), .D(count[4]), 
         .Z(n4_adj_162)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i15593_2_lut (.A(n230[3]), .B(n4), .Z(n43[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15593_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_rep_487 (.A(count[15]), .B(count[14]), .Z(n32308)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_487.init = 16'heeee;
    LUT4 i22771_2_lut_rep_428_3_lut (.A(count[15]), .B(count[14]), .C(count[12]), 
         .Z(n32249)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22771_2_lut_rep_428_3_lut.init = 16'hfefe;
    LUT4 i2_2_lut_rep_390_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(count[13]), 
         .D(count[12]), .Z(n32211)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_2_lut_rep_390_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_488 (.A(count[11]), .B(count[10]), .Z(n32309)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_488.init = 16'heeee;
    LUT4 i1_2_lut_rep_425_3_lut (.A(count[11]), .B(count[10]), .C(count[9]), 
         .Z(n32246)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_425_3_lut.init = 16'hfefe;
    LUT4 i15528_2_lut_rep_490 (.A(count[4]), .B(count[5]), .Z(n32311)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15528_2_lut_rep_490.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_272 (.A(count[4]), .B(count[5]), .C(count[7]), 
         .D(n28191), .Z(n5)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut_adj_272.init = 16'hf8f0;
    LUT4 i2_3_lut_rep_491 (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n32312)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_rep_491.init = 16'h8080;
    LUT4 i1_2_lut_rep_429_4_lut (.A(count[2]), .B(count[3]), .C(count[1]), 
         .D(count[0]), .Z(n32250)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_429_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_492 (.A(count[7]), .B(count[6]), .Z(n32313)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_492.init = 16'h8888;
    LUT4 i1_2_lut_rep_427_3_lut_4_lut (.A(count[7]), .B(count[6]), .C(count[5]), 
         .D(count[4]), .Z(n32248)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_427_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut (.A(count[7]), .B(count[6]), .C(count[5]), .Z(n29785)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i5.GSR = "ENABLED";
    LUT4 i15592_2_lut (.A(n230[2]), .B(n4), .Z(n43[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15592_2_lut.init = 16'h2222;
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i6.GSR = "ENABLED";
    LUT4 i15591_2_lut (.A(n230[1]), .B(n4), .Z(n43[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(165[10] 169[14])
    defparam i15591_2_lut.init = 16'h2222;
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n13977), .PD(n16511), .CK(debug_c_c), 
            .Q(\register[1] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam period_i0_i0.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1111), .SP(n32135), .CK(debug_c_c), .Q(n1099));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i10_3_lut_4_lut (.A(count[8]), .B(n32188), .C(n29913), .D(n29786), 
         .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i10_3_lut_4_lut.init = 16'h0100;
    IFS1P3DX latched_in_45 (.D(rc_ch1_c), .SP(n32135), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1111));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i22736_3_lut_4_lut (.A(count[8]), .B(n32188), .C(n29786), .D(n29913), 
         .Z(n30239)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i22736_3_lut_4_lut.init = 16'hfeee;
    LUT4 i1_2_lut_rep_367_3_lut_4_lut (.A(count[9]), .B(n32309), .C(n32249), 
         .D(count[13]), .Z(n32188)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_367_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut (.A(count[4]), .B(count[3]), .C(n32307), .D(n29785), 
         .Z(n29786)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfe00;
    LUT4 i22831_3_lut_4_lut (.A(n32308), .B(count[12]), .C(n32309), .D(count[13]), 
         .Z(n30334)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22831_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_273 (.A(count[0]), .B(n32312), .C(n32313), 
         .D(n32311), .Z(n29913)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_273.init = 16'h8000;
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i7.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(count[8]), .B(n32313), .C(count[5]), .D(n32247), 
         .Z(n44_adj_161)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'heaaa;
    LUT4 i23148_3_lut (.A(count[8]), .B(count[6]), .C(n5), .Z(n30318)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i23148_3_lut.init = 16'h0101;
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32135), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3AX valid_48 (.D(n32124), .SP(n28231), .CK(debug_c_c), .Q(n1105));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam valid_48.GSR = "ENABLED";
    CCU2D sub_51_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27546), 
          .S0(n230[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_9.INIT1 = 16'h0000;
    defparam sub_51_add_2_9.INJECT1_0 = "NO";
    defparam sub_51_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27545), 
          .COUT(n27546), .S0(n230[5]), .S1(n230[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_7.INJECT1_0 = "NO";
    defparam sub_51_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27544), 
          .COUT(n27545), .S0(n230[3]), .S1(n230[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_5.INJECT1_0 = "NO";
    defparam sub_51_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27543), 
          .COUT(n27544), .S0(n230[1]), .S1(n230[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_51_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_51_add_2_3.INJECT1_0 = "NO";
    defparam sub_51_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_51_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27543), 
          .S1(n230[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(168[22:33])
    defparam sub_51_add_2_1.INIT0 = 16'hF000;
    defparam sub_51_add_2_1.INIT1 = 16'h5555;
    defparam sub_51_add_2_1.INJECT1_0 = "NO";
    defparam sub_51_add_2_1.INJECT1_1 = "NO";
    CCU2D add_1763_17 (.A0(count[15]), .B0(n32274), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27114), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1763_17.INIT0 = 16'hd222;
    defparam add_1763_17.INIT1 = 16'h0000;
    defparam add_1763_17.INJECT1_0 = "NO";
    defparam add_1763_17.INJECT1_1 = "NO";
    CCU2D add_1763_15 (.A0(count[13]), .B0(n32274), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n32274), .C1(GND_net), .D1(GND_net), .CIN(n27113), 
          .COUT(n27114), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1763_15.INIT0 = 16'hd222;
    defparam add_1763_15.INIT1 = 16'hd222;
    defparam add_1763_15.INJECT1_0 = "NO";
    defparam add_1763_15.INJECT1_1 = "NO";
    CCU2D add_1763_13 (.A0(count[11]), .B0(n32274), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n32274), .C1(GND_net), .D1(GND_net), .CIN(n27112), 
          .COUT(n27113), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1763_13.INIT0 = 16'hd222;
    defparam add_1763_13.INIT1 = 16'hd222;
    defparam add_1763_13.INJECT1_0 = "NO";
    defparam add_1763_13.INJECT1_1 = "NO";
    CCU2D add_1763_11 (.A0(count[9]), .B0(n32274), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n32274), .C1(GND_net), .D1(GND_net), .CIN(n27111), 
          .COUT(n27112), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1763_11.INIT0 = 16'hd222;
    defparam add_1763_11.INIT1 = 16'hd222;
    defparam add_1763_11.INJECT1_0 = "NO";
    defparam add_1763_11.INJECT1_1 = "NO";
    CCU2D add_1763_9 (.A0(count[7]), .B0(n32274), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n32274), .C1(GND_net), .D1(GND_net), .CIN(n27110), 
          .COUT(n27111), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1763_9.INIT0 = 16'hd222;
    defparam add_1763_9.INIT1 = 16'hd222;
    defparam add_1763_9.INJECT1_0 = "NO";
    defparam add_1763_9.INJECT1_1 = "NO";
    CCU2D add_1763_7 (.A0(count[5]), .B0(n32274), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n32274), .C1(GND_net), .D1(GND_net), .CIN(n27109), 
          .COUT(n27110), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1763_7.INIT0 = 16'hd222;
    defparam add_1763_7.INIT1 = 16'hd222;
    defparam add_1763_7.INJECT1_0 = "NO";
    defparam add_1763_7.INJECT1_1 = "NO";
    CCU2D add_1763_5 (.A0(count[3]), .B0(n32274), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n32274), .C1(GND_net), .D1(GND_net), .CIN(n27108), 
          .COUT(n27109), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1763_5.INIT0 = 16'hd222;
    defparam add_1763_5.INIT1 = 16'hd222;
    defparam add_1763_5.INJECT1_0 = "NO";
    defparam add_1763_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_274 (.A(n30239), .B(n30033), .C(n32309), .D(n29667), 
         .Z(n28129)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_274.init = 16'hcecc;
    LUT4 i3_4_lut_adj_275 (.A(n54), .B(n32211), .C(n4), .D(n22550), 
         .Z(n29667)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut_adj_275.init = 16'h0010;
    LUT4 i2_4_lut_adj_276 (.A(count[13]), .B(count[12]), .C(n28276), .D(n32246), 
         .Z(n28328)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_276.init = 16'h8880;
    LUT4 i2_4_lut_adj_277 (.A(n32313), .B(count[5]), .C(count[8]), .D(n4_adj_162), 
         .Z(n28276)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_277.init = 16'ha080;
    CCU2D add_1763_3 (.A0(count[1]), .B0(n32274), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n32274), .C1(GND_net), .D1(GND_net), .CIN(n27107), 
          .COUT(n27108), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1763_3.INIT0 = 16'hd222;
    defparam add_1763_3.INIT1 = 16'hd222;
    defparam add_1763_3.INJECT1_0 = "NO";
    defparam add_1763_3.INJECT1_1 = "NO";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32135), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(137[9] 186[6])
    defparam count_i0_i3.GSR = "ENABLED";
    CCU2D add_1763_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n28288), .B1(n1111), .C1(count[0]), .D1(n1099), .COUT(n27107), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(157[7] 184[10])
    defparam add_1763_1.INIT0 = 16'hF000;
    defparam add_1763_1.INIT1 = 16'ha565;
    defparam add_1763_1.INJECT1_0 = "NO";
    defparam add_1763_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module SabertoothSerialPeripheral
//

module SabertoothSerialPeripheral (debug_c_c, n13545, n282, n32147, 
            n34066, \databus[6] , n34070, \databus[5] , \databus[4] , 
            n34067, \databus[3] , \databus[2] , \databus[1] , \databus[0] , 
            \register[0] , n13560, n32146, \read_size[0] , n2760, 
            n21718, n34068, prev_select, \select[2] , \register_addr[0] , 
            n32285, read_value, n9482, GND_net, n34065, n8447, n32227, 
            state, n29194, n11013, n34071, n29883, n107) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n13545;
    input n282;
    input n32147;
    input n34066;
    input \databus[6] ;
    input n34070;
    input \databus[5] ;
    input \databus[4] ;
    input n34067;
    input \databus[3] ;
    input \databus[2] ;
    input \databus[1] ;
    input \databus[0] ;
    output [7:0]\register[0] ;
    input n13560;
    input n32146;
    output \read_size[0] ;
    input n2760;
    input n21718;
    input n34068;
    output prev_select;
    input \select[2] ;
    input \register_addr[0] ;
    input n32285;
    output [7:0]read_value;
    input n9482;
    input GND_net;
    input n34065;
    output n8447;
    input n32227;
    output [3:0]state;
    input n29194;
    output n11013;
    input n34071;
    input n29883;
    input n107;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    wire [7:0]\register[0]_c ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(84[12:20])
    wire [7:0]n28;
    
    wire n30135, n9389;
    wire [31:0]n63;
    
    wire n32226, n28033, n9386;
    wire [7:0]n6145;
    
    FD1P3AX register_0__i16 (.D(n282), .SP(n13545), .CK(debug_c_c), .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i16.GSR = "ENABLED";
    FD1P3JX register_0__i15 (.D(\databus[6] ), .SP(n32147), .PD(n34066), 
            .CK(debug_c_c), .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i15.GSR = "ENABLED";
    FD1P3JX register_0__i14 (.D(\databus[5] ), .SP(n32147), .PD(n34070), 
            .CK(debug_c_c), .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i14.GSR = "ENABLED";
    FD1P3JX register_0__i13 (.D(\databus[4] ), .SP(n32147), .PD(n34066), 
            .CK(debug_c_c), .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i13.GSR = "ENABLED";
    FD1P3JX register_0__i12 (.D(\databus[3] ), .SP(n32147), .PD(n34067), 
            .CK(debug_c_c), .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i12.GSR = "ENABLED";
    FD1P3JX register_0__i11 (.D(\databus[2] ), .SP(n32147), .PD(n34066), 
            .CK(debug_c_c), .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i11.GSR = "ENABLED";
    FD1P3JX register_0__i10 (.D(\databus[1] ), .SP(n32147), .PD(n34067), 
            .CK(debug_c_c), .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i10.GSR = "ENABLED";
    FD1P3JX register_0__i9 (.D(\databus[0] ), .SP(n32147), .PD(n34067), 
            .CK(debug_c_c), .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i9.GSR = "ENABLED";
    FD1P3AX register_0__i8 (.D(n282), .SP(n13560), .CK(debug_c_c), .Q(\register[0] [7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i8.GSR = "ENABLED";
    FD1P3JX register_0__i7 (.D(\databus[6] ), .SP(n32146), .PD(n34067), 
            .CK(debug_c_c), .Q(\register[0]_c [6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i7.GSR = "ENABLED";
    FD1P3JX register_0__i6 (.D(\databus[5] ), .SP(n32146), .PD(n34067), 
            .CK(debug_c_c), .Q(\register[0]_c [5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i6.GSR = "ENABLED";
    FD1P3JX register_0__i5 (.D(\databus[4] ), .SP(n32146), .PD(n34067), 
            .CK(debug_c_c), .Q(\register[0]_c [4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i5.GSR = "ENABLED";
    FD1P3JX register_0__i4 (.D(\databus[3] ), .SP(n32146), .PD(n34067), 
            .CK(debug_c_c), .Q(\register[0]_c [3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i4.GSR = "ENABLED";
    FD1P3JX register_0__i3 (.D(\databus[2] ), .SP(n32146), .PD(n34067), 
            .CK(debug_c_c), .Q(\register[0]_c [2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i3.GSR = "ENABLED";
    FD1P3JX register_0__i2 (.D(\databus[1] ), .SP(n32146), .PD(n34067), 
            .CK(debug_c_c), .Q(\register[0]_c [1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i2.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n21718), .SP(n2760), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3JX register_0__i1 (.D(\databus[0] ), .SP(n32146), .PD(n34068), 
            .CK(debug_c_c), .Q(\register[0]_c [0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam register_0__i1.GSR = "ENABLED";
    FD1S3AX prev_select_138 (.D(\select[2] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam prev_select_138.GSR = "ENABLED";
    LUT4 mux_1904_Mux_1_i1_3_lut (.A(\register[0]_c [1]), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n28[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1904_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1904_Mux_2_i1_3_lut (.A(\register[0]_c [2]), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n28[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1904_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1904_Mux_3_i1_3_lut (.A(\register[0]_c [3]), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n28[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1904_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1904_Mux_4_i1_3_lut (.A(\register[0]_c [4]), .B(\register[1] [4]), 
         .C(\register_addr[0] ), .Z(n28[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1904_Mux_4_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1904_Mux_5_i1_3_lut (.A(\register[0]_c [5]), .B(\register[1] [5]), 
         .C(\register_addr[0] ), .Z(n28[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1904_Mux_5_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1904_Mux_6_i1_3_lut (.A(\register[0]_c [6]), .B(\register[1] [6]), 
         .C(\register_addr[0] ), .Z(n28[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1904_Mux_6_i1_3_lut.init = 16'hcaca;
    LUT4 i15589_4_lut_4_lut (.A(\register[1] [7]), .B(n32285), .C(n30135), 
         .D(n9389), .Z(n63[6])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(89[23:51])
    defparam i15589_4_lut_4_lut.init = 16'hffde;
    LUT4 i1_4_lut_4_lut (.A(\register[1] [7]), .B(n32285), .C(\register[1] [1]), 
         .D(n32226), .Z(n9389)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(89[23:51])
    defparam i1_4_lut_4_lut.init = 16'h2000;
    LUT4 i1_4_lut_4_lut_adj_269 (.A(\register[0] [7]), .B(n32285), .C(\register[0]_c [1]), 
         .D(n28033), .Z(n9386)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(88[22:50])
    defparam i1_4_lut_4_lut_adj_269.init = 16'h2000;
    LUT4 mux_1904_Mux_7_i1_3_lut (.A(\register[0] [7]), .B(\register[1] [7]), 
         .C(\register_addr[0] ), .Z(n6145[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1904_Mux_7_i1_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i1 (.D(n28[1]), .SP(n2760), .CD(n9482), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n28[2]), .SP(n2760), .CD(n9482), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n28[3]), .SP(n2760), .CD(n9482), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n28[4]), .SP(n2760), .CD(n9482), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n28[5]), .SP(n2760), .CD(n9482), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n28[6]), .SP(n2760), .CD(n9482), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6145[7]), .SP(n2760), .CD(n9482), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n6145[0]), .SP(n2760), .CD(n9482), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=29, LSE_RCOL=56, LSE_LLINE=530, LSE_RLINE=538 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(101[9] 139[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 mux_1904_Mux_0_i1_3_lut (.A(\register[0]_c [0]), .B(\register[1] [0]), 
         .C(\register_addr[0] ), .Z(n6145[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(112[7] 128[14])
    defparam mux_1904_Mux_0_i1_3_lut.init = 16'hcaca;
    SabertoothSerial sserial (.debug_c_c(debug_c_c), .GND_net(GND_net), 
            .n89(n63[6]), .\register[1][2] (\register[1] [2]), .\register[1][1] (\register[1] [1]), 
            .\register[1][4] (\register[1] [4]), .\register[1][3] (\register[1] [3]), 
            .\register[0][2] (\register[0]_c [2]), .\register[0][1] (\register[0]_c [1]), 
            .\register[0][3] (\register[0]_c [3]), .\register[0][4] (\register[0]_c [4]), 
            .\register[0][7] (\register[0] [7]), .n34065(n34065), .n8447(n8447), 
            .n9389(n9389), .n32285(n32285), .n9386(n9386), .\register[1][5] (\register[1] [5]), 
            .\register[1][6] (\register[1] [6]), .n32226(n32226), .\register[1][7] (\register[1] [7]), 
            .\register[0][5] (\register[0]_c [5]), .n30135(n30135), .\register[0][6] (\register[0]_c [6]), 
            .n32227(n32227), .n28033(n28033), .state({state}), .n34066(n34066), 
            .n29194(n29194), .n11013(n11013), .n34071(n34071), .n29883(n29883), 
            .n107(n107)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(142[19] 147[34])
    
endmodule
//
// Verilog Description of module SabertoothSerial
//

module SabertoothSerial (debug_c_c, GND_net, n89, \register[1][2] , 
            \register[1][1] , \register[1][4] , \register[1][3] , \register[0][2] , 
            \register[0][1] , \register[0][3] , \register[0][4] , \register[0][7] , 
            n34065, n8447, n9389, n32285, n9386, \register[1][5] , 
            \register[1][6] , n32226, \register[1][7] , \register[0][5] , 
            n30135, \register[0][6] , n32227, n28033, state, n34066, 
            n29194, n11013, n34071, n29883, n107) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input GND_net;
    input n89;
    input \register[1][2] ;
    input \register[1][1] ;
    input \register[1][4] ;
    input \register[1][3] ;
    input \register[0][2] ;
    input \register[0][1] ;
    input \register[0][3] ;
    input \register[0][4] ;
    input \register[0][7] ;
    input n34065;
    output n8447;
    input n9389;
    input n32285;
    input n9386;
    input \register[1][5] ;
    input \register[1][6] ;
    output n32226;
    input \register[1][7] ;
    input \register[0][5] ;
    output n30135;
    input \register[0][6] ;
    input n32227;
    output n28033;
    output [3:0]state;
    input n34066;
    input n29194;
    output n11013;
    input n34071;
    input n29883;
    input n107;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n1096, n32136, n32277;
    wire [7:0]n5445;
    
    wire n7;
    wire [7:0]n5454;
    
    wire n29636, n6, n28970;
    wire [31:0]n63;
    wire [3:0]state_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(17[12:17])
    wire [3:0]n16;
    
    wire n32272, n32197, n32225, n32273, n32228, n11343, n32198, 
        n12191, n12_adj_156, n32171, select_clk, n14170, n11889, 
        n32170, n29563, n20, n12329, n11260;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(16[12:19])
    
    wire n32128, n12327;
    wire [3:0]n7749;
    
    wire n24, n10193, n6_adj_157, n29565;
    
    FD1P3IX send_31 (.D(n32277), .SP(n32136), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1096));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam send_31.GSR = "ENABLED";
    PFUMX mux_1837_i7 (.BLUT(n89), .ALUT(n5445[6]), .C0(n7), .Z(n5454[6]));
    PFUMX i30 (.BLUT(n29636), .ALUT(n6), .C0(n7), .Z(n28970));
    PFUMX mux_1837_i2 (.BLUT(n63[1]), .ALUT(n5445[1]), .C0(n7), .Z(n5454[1]));
    FD1S3IX state__i0 (.D(n16[0]), .CK(debug_c_c), .CD(GND_net), .Q(state_c[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam state__i0.GSR = "ENABLED";
    PFUMX mux_1837_i3 (.BLUT(n63[2]), .ALUT(n5445[2]), .C0(n7), .Z(n5454[2]));
    PFUMX mux_1837_i4 (.BLUT(n63[3]), .ALUT(n5445[3]), .C0(n7), .Z(n5454[3]));
    PFUMX mux_1837_i5 (.BLUT(n63[4]), .ALUT(n5445[4]), .C0(n7), .Z(n5454[4]));
    PFUMX mux_1837_i6 (.BLUT(n63[5]), .ALUT(n5445[5]), .C0(n7), .Z(n5454[5]));
    LUT4 i4383_2_lut_rep_451 (.A(\register[1][2] ), .B(\register[1][1] ), 
         .Z(n32272)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4383_2_lut_rep_451.init = 16'h8888;
    LUT4 i5439_2_lut_rep_376_3_lut_4_lut (.A(\register[1][2] ), .B(\register[1][1] ), 
         .C(\register[1][4] ), .D(\register[1][3] ), .Z(n32197)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5439_2_lut_rep_376_3_lut_4_lut.init = 16'h8000;
    LUT4 i4390_2_lut_rep_404_3_lut (.A(\register[1][2] ), .B(\register[1][1] ), 
         .C(\register[1][3] ), .Z(n32225)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i4390_2_lut_rep_404_3_lut.init = 16'h8080;
    LUT4 i4598_2_lut_rep_452 (.A(\register[0][2] ), .B(\register[0][1] ), 
         .Z(n32273)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4598_2_lut_rep_452.init = 16'h8888;
    LUT4 i4618_2_lut_rep_407_3_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][3] ), .Z(n32228)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i4618_2_lut_rep_407_3_lut.init = 16'h8080;
    LUT4 i4626_2_lut_3_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][3] ), .Z(n11343)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i4626_2_lut_3_lut.init = 16'h7878;
    LUT4 i5592_2_lut_rep_377_3_lut_4_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][4] ), .D(\register[0][3] ), .Z(n32198)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5592_2_lut_rep_377_3_lut_4_lut.init = 16'h8000;
    LUT4 i5471_2_lut_3_lut_4_lut (.A(\register[0][2] ), .B(\register[0][1] ), 
         .C(\register[0][4] ), .D(\register[0][3] ), .Z(n12191)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i5471_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i4059_1_lut_rep_456 (.A(state_c[0]), .Z(n32277)) /* synthesis lut_function=(!(A)) */ ;
    defparam i4059_1_lut_rep_456.init = 16'h5555;
    LUT4 i6_4_lut_4_lut (.A(state_c[0]), .B(\register[0][7] ), .C(n12_adj_156), 
         .D(n32171), .Z(n6)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i6_4_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_4_lut_4_lut (.A(state_c[0]), .B(select_clk), .C(n34065), 
         .D(n8447), .Z(n14170)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut_4_lut.init = 16'h0100;
    LUT4 i15585_4_lut (.A(\register[1][3] ), .B(n9389), .C(n32285), .D(n32272), 
         .Z(n63[2])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15585_4_lut.init = 16'hcdce;
    LUT4 i15106_4_lut (.A(n11343), .B(n11889), .C(n9386), .D(n32285), 
         .Z(n5445[2])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i15106_4_lut.init = 16'h3032;
    LUT4 i5452_2_lut_rep_349_3_lut_4_lut (.A(\register[1][3] ), .B(n32272), 
         .C(\register[1][5] ), .D(\register[1][4] ), .Z(n32170)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5452_2_lut_rep_349_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_405 (.A(\register[1][6] ), .B(n29563), .Z(n32226)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_405.init = 16'h8888;
    LUT4 i1_3_lut_4_lut (.A(\register[1][6] ), .B(n29563), .C(\register[1][7] ), 
         .D(\register[1][1] ), .Z(n20)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h80ff;
    LUT4 i5594_2_lut_rep_350_3_lut_4_lut (.A(\register[0][3] ), .B(n32273), 
         .C(\register[0][5] ), .D(\register[0][4] ), .Z(n32171)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5594_2_lut_rep_350_3_lut_4_lut.init = 16'h8000;
    LUT4 i5609_2_lut_3_lut_4_lut (.A(\register[0][3] ), .B(n32273), .C(\register[0][5] ), 
         .D(\register[0][4] ), .Z(n12329)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i5609_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i15584_4_lut (.A(\register[1][2] ), .B(n9389), .C(n32285), .D(\register[1][1] ), 
         .Z(n63[1])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15584_4_lut.init = 16'hcdce;
    LUT4 i15105_4_lut (.A(n11260), .B(n11889), .C(n9386), .D(n32285), 
         .Z(n5445[1])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i15105_4_lut.init = 16'h3032;
    LUT4 i4543_2_lut (.A(\register[0][2] ), .B(\register[0][1] ), .Z(n11260)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4543_2_lut.init = 16'h6666;
    FD1P3AX tx_data_i0_i0 (.D(n32128), .SP(n14170), .CK(debug_c_c), .Q(tx_data[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    LUT4 i15586_4_lut (.A(\register[1][4] ), .B(n9389), .C(n32285), .D(n32225), 
         .Z(n63[3])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15586_4_lut.init = 16'hcdce;
    LUT4 i15107_4_lut (.A(n12191), .B(n11889), .C(n9386), .D(n32285), 
         .Z(n5445[3])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i15107_4_lut.init = 16'h3032;
    LUT4 i15587_4_lut (.A(\register[1][5] ), .B(n9389), .C(n32285), .D(n32197), 
         .Z(n63[4])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15587_4_lut.init = 16'hcdce;
    LUT4 i15108_4_lut (.A(n12329), .B(n11889), .C(n9386), .D(n32285), 
         .Z(n5445[4])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i15108_4_lut.init = 16'h3032;
    LUT4 i15588_4_lut (.A(\register[1][6] ), .B(n9389), .C(n32285), .D(n32170), 
         .Z(n63[5])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(48[20:75])
    defparam i15588_4_lut.init = 16'hcdce;
    LUT4 i22639_2_lut_3_lut_4_lut (.A(\register[1][4] ), .B(n32225), .C(\register[1][6] ), 
         .D(\register[1][5] ), .Z(n30135)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22639_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i15109_4_lut (.A(n12327), .B(n11889), .C(n9386), .D(n32285), 
         .Z(n5445[5])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i15109_4_lut.init = 16'h3032;
    LUT4 i5607_2_lut_3_lut_4_lut (.A(\register[0][4] ), .B(n32228), .C(\register[0][6] ), 
         .D(\register[0][5] ), .Z(n12327)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i5607_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1P3IX state__i1 (.D(n7749[1]), .SP(n32136), .CD(GND_net), .CK(debug_c_c), 
            .Q(state_c[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam state__i1.GSR = "ENABLED";
    LUT4 n20_bdd_4_lut (.A(n20), .B(n24), .C(n7), .D(n32285), .Z(n32128)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n20_bdd_4_lut.init = 16'h00ca;
    LUT4 i4366_2_lut (.A(state_c[0]), .B(state_c[1]), .Z(n7749[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(34[6] 57[13])
    defparam i4366_2_lut.init = 16'h6666;
    FD1P3AX tx_data_i0_i1 (.D(n5454[1]), .SP(n14170), .CK(debug_c_c), 
            .Q(tx_data[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    LUT4 i15110_4_lut (.A(n32227), .B(n11889), .C(n9386), .D(n10193), 
         .Z(n5445[6])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C+(D))))) */ ;
    defparam i15110_4_lut.init = 16'h3132;
    LUT4 equal_16_i5_2_lut (.A(state_c[0]), .B(state_c[1]), .Z(n7)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(46[7:11])
    defparam equal_16_i5_2_lut.init = 16'hbbbb;
    FD1P3AX tx_data_i0_i2 (.D(n5454[2]), .SP(n14170), .CK(debug_c_c), 
            .Q(tx_data[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n5454[3]), .SP(n14170), .CK(debug_c_c), 
            .Q(tx_data[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i4 (.D(n5454[4]), .SP(n14170), .CK(debug_c_c), 
            .Q(tx_data[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i5 (.D(n5454[5]), .SP(n14170), .CK(debug_c_c), 
            .Q(tx_data[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i6 (.D(n5454[6]), .SP(n14170), .CK(debug_c_c), 
            .Q(tx_data[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i7 (.D(n28970), .SP(n14170), .CK(debug_c_c), .Q(tx_data[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n11889), .B(\register[0][1] ), .C(n28033), .D(\register[0][7] ), 
         .Z(n24)) /* synthesis lut_function=(!(A+!((C (D))+!B))) */ ;
    defparam i1_4_lut.init = 16'h5111;
    LUT4 i4385_2_lut (.A(state_c[0]), .B(state_c[1]), .Z(n11889)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i4385_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_rep_315 (.A(n8447), .B(n34065), .C(select_clk), .Z(n32136)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i2_3_lut_rep_315.init = 16'h0202;
    LUT4 i5612_2_lut_4_lut (.A(n8447), .B(n34065), .C(select_clk), .D(state_c[0]), 
         .Z(n16[0])) /* synthesis lut_function=(A (B (D)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(25[9] 61[6])
    defparam i5612_2_lut_4_lut.init = 16'hfd02;
    LUT4 i15814_3_lut_4_lut (.A(\register[0][5] ), .B(n32198), .C(n32285), 
         .D(\register[0][6] ), .Z(n10193)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i15814_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i3_4_lut (.A(\register[1][5] ), .B(\register[1][3] ), .C(\register[1][4] ), 
         .D(\register[1][2] ), .Z(n29563)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i4_4_lut (.A(\register[0][4] ), .B(\register[0][2] ), .C(\register[0][3] ), 
         .D(n6_adj_157), .Z(n28033)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i4_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_267 (.A(n32285), .B(\register[1][7] ), .C(n30135), 
         .D(n29565), .Z(n29636)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_267.init = 16'hffbf;
    LUT4 i1_2_lut (.A(\register[0][5] ), .B(\register[0][6] ), .Z(n6_adj_157)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_268 (.A(\register[1][1] ), .B(n29563), .Z(n29565)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_268.init = 16'h8888;
    LUT4 i5_4_lut (.A(\register[0][6] ), .B(state_c[1]), .C(n9386), .D(n32285), 
         .Z(n12_adj_156)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i5_4_lut.init = 16'h0002;
    \UARTTransmitter(baud_div=1250)  sender (.state({state}), .n34066(n34066), 
            .n29194(n29194), .tx_data({tx_data}), .n1096(n1096), .n34065(n34065), 
            .n11013(n11013), .n34071(n34071), .n29883(n29883), .debug_c_c(debug_c_c), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(63[26] 67[47])
    \ClockDividerP(factor=12000)  baud_gen (.select_clk(select_clk), .debug_c_c(debug_c_c), 
            .n107(n107), .GND_net(GND_net), .n8447(n8447), .n34065(n34065)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/motor-serial.v(21[25] 23[48])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=1250) 
//

module \UARTTransmitter(baud_div=1250)  (state, n34066, n29194, tx_data, 
            n1096, n34065, n11013, n34071, n29883, debug_c_c, GND_net) /* synthesis syn_module_defined=1 */ ;
    output [3:0]state;
    input n34066;
    input n29194;
    input [7:0]tx_data;
    input n1096;
    input n34065;
    output n11013;
    input n34071;
    input n29883;
    input debug_c_c;
    input GND_net;
    
    wire bclk /* synthesis SET_AS_NETWORK=\motor_serial/sserial/sender/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n31573, n31572, n31574, n31865, n13615;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n9393, n19804, n30405, n30406, n30407, n4, n27859, n5, 
        n7, n33, n19792, n34, n19798, n10, n29664;
    wire [3:0]n11;
    
    wire n12;
    
    PFUMX i23451 (.BLUT(n31573), .ALUT(n31572), .C0(state[2]), .Z(n31574));
    FD1S3IX state__i0 (.D(n31574), .CK(bclk), .CD(n34066), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    LUT4 state_1__bdd_4_lut (.A(state[1]), .B(state[0]), .C(state[3]), 
         .D(state[2]), .Z(n31865)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C (D))+!B (C (D)+!C !(D))))) */ ;
    defparam state_1__bdd_4_lut.init = 16'h0f7e;
    FD1P3AX state__i3 (.D(n29194), .SP(n13615), .CK(bclk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n9393), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut (.A(state[1]), .B(state[3]), .C(n1096), .Z(n19804)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    PFUMX i22904 (.BLUT(n30405), .ALUT(n30406), .C0(state[0]), .Z(n30407));
    LUT4 i2_4_lut (.A(n19804), .B(n4), .C(n27859), .D(state[0]), .Z(n13615)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B+!(C+!(D)))) */ ;
    defparam i2_4_lut.init = 16'hcfee;
    LUT4 i1_2_lut (.A(state[2]), .B(n34065), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i2_3_lut (.A(state[1]), .B(n1096), .C(state[3]), .Z(n27859)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i22902_4_lut (.A(n5), .B(state[1]), .C(state[3]), .D(tdata[6]), 
         .Z(n30405)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i22902_4_lut.init = 16'hfaca;
    LUT4 i22903_4_lut (.A(n7), .B(state[1]), .C(state[3]), .D(tdata[7]), 
         .Z(n30406)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i22903_4_lut.init = 16'hfaca;
    LUT4 state_1__bdd_4_lut_23596 (.A(state[1]), .B(state[0]), .C(state[3]), 
         .D(n1096), .Z(n31573)) /* synthesis lut_function=(A ((C (D))+!B)+!A !(B+!(C+(D)))) */ ;
    defparam state_1__bdd_4_lut_23596.init = 16'hb332;
    FD1P3JX tx_35 (.D(n30407), .SP(n31865), .PD(n34071), .CK(bclk), 
            .Q(n11013)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_264 (.A(state[1]), .B(tdata[0]), .Z(n33)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i1_2_lut_adj_264.init = 16'h8888;
    LUT4 i13085_3_lut (.A(tdata[2]), .B(tdata[4]), .C(state[1]), .Z(n19792)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    defparam i13085_3_lut.init = 16'hcaca;
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n9393), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n9393), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n9393), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n9393), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n9393), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n9393), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n9393), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_265 (.A(state[1]), .B(tdata[1]), .Z(n34)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i1_2_lut_adj_265.init = 16'h8888;
    LUT4 i13091_3_lut (.A(tdata[3]), .B(tdata[5]), .C(state[1]), .Z(n19798)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    defparam i13091_3_lut.init = 16'hcaca;
    LUT4 i5_3_lut (.A(state[3]), .B(n10), .C(n34065), .Z(n9393)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i5_3_lut.init = 16'h0404;
    LUT4 i4_4_lut (.A(state[2]), .B(n1096), .C(state[0]), .D(state[1]), 
         .Z(n10)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i4_4_lut.init = 16'h0004;
    FD1P3AX state__i1 (.D(n29664), .SP(n13615), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    FD1P3AX state__i2 (.D(n11[2]), .SP(n13615), .CK(bclk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=26, LSE_RCOL=47, LSE_LLINE=63, LSE_RLINE=67 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n34065), .B(state[2]), .C(n12), .D(state[3]), 
         .Z(n29664)) /* synthesis lut_function=(!(A+(B ((D)+!C)+!B !(C)))) */ ;
    defparam i1_4_lut.init = 16'h1050;
    LUT4 i22_2_lut (.A(state[1]), .B(state[0]), .Z(n12)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i22_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_266 (.A(n34065), .B(n29883), .C(state[3]), .D(state[2]), 
         .Z(n11[2])) /* synthesis lut_function=(!(A+(B (D)+!B (C+!(D))))) */ ;
    defparam i1_4_lut_adj_266.init = 16'h0144;
    LUT4 state_1__bdd_2_lut (.A(state[0]), .B(state[3]), .Z(n31572)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_1__bdd_2_lut.init = 16'h1111;
    PFUMX i5 (.BLUT(n33), .ALUT(n19792), .C0(state[2]), .Z(n5));
    PFUMX i7 (.BLUT(n34), .ALUT(n19798), .C0(state[2]), .Z(n7));
    \ClockDividerP(factor=1250)  baud_gen (.bclk(bclk), .debug_c_c(debug_c_c), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=1250) 
//

module \ClockDividerP(factor=1250)  (bclk, debug_c_c, GND_net) /* synthesis syn_module_defined=1 */ ;
    output bclk;
    input debug_c_c;
    input GND_net;
    
    wire bclk /* synthesis SET_AS_NETWORK=\motor_serial/sserial/sender/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n8482, n27780;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n27779, n27778, n27777, n27776, n27775, n27774, n27773, 
        n27772, n27771, n27770, n27769, n27768, n27767, n27766, 
        n27726;
    wire [31:0]n102;
    
    wire n27725, n27724, n27723, n27722, n27721, n27720, n27719, 
        n16571, n27718, n27717, n27716, n27715, n27714, n27713, 
        n27712, n27711, n28408, n8, n39, n52, n48, n40, n31, 
        n50, n44, n32, n42, n46, n36;
    
    FD1S3AX clk_o_14 (.D(n8482), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D add_20291_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27780), 
          .S1(n8482));
    defparam add_20291_32.INIT0 = 16'h5555;
    defparam add_20291_32.INIT1 = 16'h0000;
    defparam add_20291_32.INJECT1_0 = "NO";
    defparam add_20291_32.INJECT1_1 = "NO";
    CCU2D add_20291_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27779), .COUT(n27780));
    defparam add_20291_30.INIT0 = 16'h5555;
    defparam add_20291_30.INIT1 = 16'h5555;
    defparam add_20291_30.INJECT1_0 = "NO";
    defparam add_20291_30.INJECT1_1 = "NO";
    CCU2D add_20291_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27778), .COUT(n27779));
    defparam add_20291_28.INIT0 = 16'h5555;
    defparam add_20291_28.INIT1 = 16'h5555;
    defparam add_20291_28.INJECT1_0 = "NO";
    defparam add_20291_28.INJECT1_1 = "NO";
    CCU2D add_20291_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27777), .COUT(n27778));
    defparam add_20291_26.INIT0 = 16'h5555;
    defparam add_20291_26.INIT1 = 16'h5555;
    defparam add_20291_26.INJECT1_0 = "NO";
    defparam add_20291_26.INJECT1_1 = "NO";
    CCU2D add_20291_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27776), .COUT(n27777));
    defparam add_20291_24.INIT0 = 16'h5555;
    defparam add_20291_24.INIT1 = 16'h5555;
    defparam add_20291_24.INJECT1_0 = "NO";
    defparam add_20291_24.INJECT1_1 = "NO";
    CCU2D add_20291_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27775), .COUT(n27776));
    defparam add_20291_22.INIT0 = 16'h5555;
    defparam add_20291_22.INIT1 = 16'h5555;
    defparam add_20291_22.INJECT1_0 = "NO";
    defparam add_20291_22.INJECT1_1 = "NO";
    CCU2D add_20291_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27774), .COUT(n27775));
    defparam add_20291_20.INIT0 = 16'h5555;
    defparam add_20291_20.INIT1 = 16'h5555;
    defparam add_20291_20.INJECT1_0 = "NO";
    defparam add_20291_20.INJECT1_1 = "NO";
    CCU2D add_20291_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27773), .COUT(n27774));
    defparam add_20291_18.INIT0 = 16'h5555;
    defparam add_20291_18.INIT1 = 16'h5555;
    defparam add_20291_18.INJECT1_0 = "NO";
    defparam add_20291_18.INJECT1_1 = "NO";
    CCU2D add_20291_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27772), .COUT(n27773));
    defparam add_20291_16.INIT0 = 16'h5555;
    defparam add_20291_16.INIT1 = 16'h5555;
    defparam add_20291_16.INJECT1_0 = "NO";
    defparam add_20291_16.INJECT1_1 = "NO";
    CCU2D add_20291_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27771), .COUT(n27772));
    defparam add_20291_14.INIT0 = 16'h5555;
    defparam add_20291_14.INIT1 = 16'h5555;
    defparam add_20291_14.INJECT1_0 = "NO";
    defparam add_20291_14.INJECT1_1 = "NO";
    CCU2D add_20291_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27770), .COUT(n27771));
    defparam add_20291_12.INIT0 = 16'h5555;
    defparam add_20291_12.INIT1 = 16'h5555;
    defparam add_20291_12.INJECT1_0 = "NO";
    defparam add_20291_12.INJECT1_1 = "NO";
    CCU2D add_20291_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27769), .COUT(n27770));
    defparam add_20291_10.INIT0 = 16'h5aaa;
    defparam add_20291_10.INIT1 = 16'h5555;
    defparam add_20291_10.INJECT1_0 = "NO";
    defparam add_20291_10.INJECT1_1 = "NO";
    CCU2D add_20291_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27768), 
          .COUT(n27769));
    defparam add_20291_8.INIT0 = 16'h5555;
    defparam add_20291_8.INIT1 = 16'h5555;
    defparam add_20291_8.INJECT1_0 = "NO";
    defparam add_20291_8.INJECT1_1 = "NO";
    CCU2D add_20291_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27767), 
          .COUT(n27768));
    defparam add_20291_6.INIT0 = 16'h5aaa;
    defparam add_20291_6.INIT1 = 16'h5aaa;
    defparam add_20291_6.INJECT1_0 = "NO";
    defparam add_20291_6.INJECT1_1 = "NO";
    CCU2D add_20291_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27766), 
          .COUT(n27767));
    defparam add_20291_4.INIT0 = 16'h5555;
    defparam add_20291_4.INIT1 = 16'h5aaa;
    defparam add_20291_4.INJECT1_0 = "NO";
    defparam add_20291_4.INJECT1_1 = "NO";
    CCU2D add_20291_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27766));
    defparam add_20291_2.INIT0 = 16'h1000;
    defparam add_20291_2.INIT1 = 16'h5555;
    defparam add_20291_2.INJECT1_0 = "NO";
    defparam add_20291_2.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27726), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_33.INIT1 = 16'h0000;
    defparam count_2669_add_4_33.INJECT1_0 = "NO";
    defparam count_2669_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27725), .COUT(n27726), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2669_add_4_31.INJECT1_0 = "NO";
    defparam count_2669_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27724), .COUT(n27725), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2669_add_4_29.INJECT1_0 = "NO";
    defparam count_2669_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27723), .COUT(n27724), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2669_add_4_27.INJECT1_0 = "NO";
    defparam count_2669_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27722), .COUT(n27723), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2669_add_4_25.INJECT1_0 = "NO";
    defparam count_2669_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27721), .COUT(n27722), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2669_add_4_23.INJECT1_0 = "NO";
    defparam count_2669_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27720), .COUT(n27721), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2669_add_4_21.INJECT1_0 = "NO";
    defparam count_2669_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27719), .COUT(n27720), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2669_add_4_19.INJECT1_0 = "NO";
    defparam count_2669_add_4_19.INJECT1_1 = "NO";
    FD1S3IX count_2669__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i0.GSR = "ENABLED";
    CCU2D count_2669_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27718), .COUT(n27719), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2669_add_4_17.INJECT1_0 = "NO";
    defparam count_2669_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27717), .COUT(n27718), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2669_add_4_15.INJECT1_0 = "NO";
    defparam count_2669_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27716), .COUT(n27717), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2669_add_4_13.INJECT1_0 = "NO";
    defparam count_2669_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27715), .COUT(n27716), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2669_add_4_11.INJECT1_0 = "NO";
    defparam count_2669_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27714), .COUT(n27715), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2669_add_4_9.INJECT1_0 = "NO";
    defparam count_2669_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27713), .COUT(n27714), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2669_add_4_7.INJECT1_0 = "NO";
    defparam count_2669_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27712), .COUT(n27713), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2669_add_4_5.INJECT1_0 = "NO";
    defparam count_2669_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27711), .COUT(n27712), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2669_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2669_add_4_3.INJECT1_0 = "NO";
    defparam count_2669_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2669_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27711), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669_add_4_1.INIT0 = 16'hF000;
    defparam count_2669_add_4_1.INIT1 = 16'h0555;
    defparam count_2669_add_4_1.INJECT1_0 = "NO";
    defparam count_2669_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2669__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i1.GSR = "ENABLED";
    LUT4 i23128_4_lut (.A(n28408), .B(count[5]), .C(n8), .D(count[0]), 
         .Z(n16571)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23128_4_lut.init = 16'h4000;
    LUT4 i26_4_lut (.A(n39), .B(n52), .C(n48), .D(n40), .Z(n28408)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i3_3_lut (.A(count[10]), .B(count[6]), .C(count[7]), .Z(n8)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i3_3_lut.init = 16'h8080;
    LUT4 i12_2_lut (.A(count[30]), .B(count[13]), .Z(n39)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i12_2_lut.init = 16'heeee;
    LUT4 i25_4_lut (.A(n31), .B(n50), .C(n44), .D(n32), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(count[27]), .B(n42), .C(count[23]), .D(count[17]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(count[22]), .B(count[18]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i4_2_lut (.A(count[28]), .B(count[9]), .Z(n31)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(count[19]), .B(n46), .C(n36), .D(count[25]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(count[4]), .B(count[11]), .C(count[8]), .D(count[14]), 
         .Z(n44)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(count[12]), .B(count[1]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i19_4_lut (.A(count[20]), .B(count[2]), .C(count[24]), .D(count[29]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(count[26]), .B(count[3]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i15_4_lut (.A(count[16]), .B(count[15]), .C(count[31]), .D(count[21]), 
         .Z(n42)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i15_4_lut.init = 16'hfffe;
    FD1S3IX count_2669__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i2.GSR = "ENABLED";
    FD1S3IX count_2669__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i3.GSR = "ENABLED";
    FD1S3IX count_2669__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i4.GSR = "ENABLED";
    FD1S3IX count_2669__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i5.GSR = "ENABLED";
    FD1S3IX count_2669__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i6.GSR = "ENABLED";
    FD1S3IX count_2669__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i7.GSR = "ENABLED";
    FD1S3IX count_2669__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i8.GSR = "ENABLED";
    FD1S3IX count_2669__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i9.GSR = "ENABLED";
    FD1S3IX count_2669__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i10.GSR = "ENABLED";
    FD1S3IX count_2669__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i11.GSR = "ENABLED";
    FD1S3IX count_2669__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i12.GSR = "ENABLED";
    FD1S3IX count_2669__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i13.GSR = "ENABLED";
    FD1S3IX count_2669__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i14.GSR = "ENABLED";
    FD1S3IX count_2669__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i15.GSR = "ENABLED";
    FD1S3IX count_2669__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i16.GSR = "ENABLED";
    FD1S3IX count_2669__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i17.GSR = "ENABLED";
    FD1S3IX count_2669__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i18.GSR = "ENABLED";
    FD1S3IX count_2669__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i19.GSR = "ENABLED";
    FD1S3IX count_2669__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i20.GSR = "ENABLED";
    FD1S3IX count_2669__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i21.GSR = "ENABLED";
    FD1S3IX count_2669__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i22.GSR = "ENABLED";
    FD1S3IX count_2669__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i23.GSR = "ENABLED";
    FD1S3IX count_2669__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i24.GSR = "ENABLED";
    FD1S3IX count_2669__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i25.GSR = "ENABLED";
    FD1S3IX count_2669__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i26.GSR = "ENABLED";
    FD1S3IX count_2669__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i27.GSR = "ENABLED";
    FD1S3IX count_2669__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i28.GSR = "ENABLED";
    FD1S3IX count_2669__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i29.GSR = "ENABLED";
    FD1S3IX count_2669__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i30.GSR = "ENABLED";
    FD1S3IX count_2669__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n16571), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2669__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000) 
//

module \ClockDividerP(factor=12000)  (select_clk, debug_c_c, n107, GND_net, 
            n8447, n34065) /* synthesis syn_module_defined=1 */ ;
    output select_clk;
    input debug_c_c;
    input n107;
    input GND_net;
    output n8447;
    input n34065;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n40, n34, n30336, n42, n38, n30, n36, n26, n30250, 
        n2907;
    wire [31:0]n134;
    
    wire n27765, n27764, n27763, n27762, n27761, n27760, n27759, 
        n27758, n27757, n27756, n27755, n27754, n30446, n29640, 
        n30186, n29, n27753, n27710, n27709, n27708, n27707, n27706, 
        n27705, n27704, n27703, n27702, n27701, n27700, n27699, 
        n27698, n27697, n27696, n27695;
    
    LUT4 i20_4_lut (.A(count[31]), .B(n40), .C(n34), .D(n30336), .Z(n42)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i20_4_lut.init = 16'hfeff;
    LUT4 i16_4_lut (.A(count[20]), .B(count[23]), .C(count[15]), .D(count[29]), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(count[22]), .B(count[5]), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i18_4_lut (.A(count[21]), .B(n36), .C(n26), .D(count[25]), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i12_4_lut (.A(count[28]), .B(count[8]), .C(count[18]), .D(count[16]), 
         .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i22833_4_lut (.A(count[10]), .B(count[3]), .C(count[13]), .D(n30250), 
         .Z(n30336)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22833_4_lut.init = 16'h8000;
    LUT4 i22747_2_lut (.A(count[0]), .B(count[4]), .Z(n30250)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22747_2_lut.init = 16'h8888;
    LUT4 i14_4_lut (.A(count[17]), .B(count[27]), .C(count[24]), .D(count[30]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(count[26]), .B(count[12]), .Z(n26)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i4_2_lut.init = 16'heeee;
    FD1S3AX clk_o_14 (.D(n107), .CK(debug_c_c), .Q(select_clk)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=25, LSE_RCOL=48, LSE_LLINE=21, LSE_RLINE=23 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2668__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2907), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i0.GSR = "ENABLED";
    CCU2D add_20292_28 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27765), 
          .S1(n8447));
    defparam add_20292_28.INIT0 = 16'h5555;
    defparam add_20292_28.INIT1 = 16'h0000;
    defparam add_20292_28.INJECT1_0 = "NO";
    defparam add_20292_28.INJECT1_1 = "NO";
    CCU2D add_20292_26 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27764), .COUT(n27765));
    defparam add_20292_26.INIT0 = 16'h5555;
    defparam add_20292_26.INIT1 = 16'h5555;
    defparam add_20292_26.INJECT1_0 = "NO";
    defparam add_20292_26.INJECT1_1 = "NO";
    CCU2D add_20292_24 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27763), .COUT(n27764));
    defparam add_20292_24.INIT0 = 16'h5555;
    defparam add_20292_24.INIT1 = 16'h5555;
    defparam add_20292_24.INJECT1_0 = "NO";
    defparam add_20292_24.INJECT1_1 = "NO";
    CCU2D add_20292_22 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27762), .COUT(n27763));
    defparam add_20292_22.INIT0 = 16'h5555;
    defparam add_20292_22.INIT1 = 16'h5555;
    defparam add_20292_22.INJECT1_0 = "NO";
    defparam add_20292_22.INJECT1_1 = "NO";
    CCU2D add_20292_20 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27761), .COUT(n27762));
    defparam add_20292_20.INIT0 = 16'h5555;
    defparam add_20292_20.INIT1 = 16'h5555;
    defparam add_20292_20.INJECT1_0 = "NO";
    defparam add_20292_20.INJECT1_1 = "NO";
    CCU2D add_20292_18 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27760), .COUT(n27761));
    defparam add_20292_18.INIT0 = 16'h5555;
    defparam add_20292_18.INIT1 = 16'h5555;
    defparam add_20292_18.INJECT1_0 = "NO";
    defparam add_20292_18.INJECT1_1 = "NO";
    CCU2D add_20292_16 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27759), .COUT(n27760));
    defparam add_20292_16.INIT0 = 16'h5555;
    defparam add_20292_16.INIT1 = 16'h5555;
    defparam add_20292_16.INJECT1_0 = "NO";
    defparam add_20292_16.INJECT1_1 = "NO";
    CCU2D add_20292_14 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27758), .COUT(n27759));
    defparam add_20292_14.INIT0 = 16'h5555;
    defparam add_20292_14.INIT1 = 16'h5555;
    defparam add_20292_14.INJECT1_0 = "NO";
    defparam add_20292_14.INJECT1_1 = "NO";
    CCU2D add_20292_12 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27757), .COUT(n27758));
    defparam add_20292_12.INIT0 = 16'h5555;
    defparam add_20292_12.INIT1 = 16'h5555;
    defparam add_20292_12.INJECT1_0 = "NO";
    defparam add_20292_12.INJECT1_1 = "NO";
    CCU2D add_20292_10 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27756), .COUT(n27757));
    defparam add_20292_10.INIT0 = 16'h5555;
    defparam add_20292_10.INIT1 = 16'h5555;
    defparam add_20292_10.INJECT1_0 = "NO";
    defparam add_20292_10.INJECT1_1 = "NO";
    CCU2D add_20292_8 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27755), .COUT(n27756));
    defparam add_20292_8.INIT0 = 16'h5555;
    defparam add_20292_8.INIT1 = 16'h5aaa;
    defparam add_20292_8.INJECT1_0 = "NO";
    defparam add_20292_8.INJECT1_1 = "NO";
    CCU2D add_20292_6 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27754), .COUT(n27755));
    defparam add_20292_6.INIT0 = 16'h5aaa;
    defparam add_20292_6.INIT1 = 16'h5aaa;
    defparam add_20292_6.INJECT1_0 = "NO";
    defparam add_20292_6.INJECT1_1 = "NO";
    LUT4 i23046_2_lut (.A(n30446), .B(n34065), .Z(n2907)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23046_2_lut.init = 16'heeee;
    LUT4 i23044_4_lut (.A(n29640), .B(count[9]), .C(n30186), .D(count[6]), 
         .Z(n30446)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i23044_4_lut.init = 16'h4000;
    LUT4 i21_4_lut (.A(n29), .B(n42), .C(n38), .D(n30), .Z(n29640)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i22688_4_lut (.A(count[2]), .B(count[11]), .C(count[1]), .D(count[7]), 
         .Z(n30186)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22688_4_lut.init = 16'h8000;
    LUT4 i7_2_lut (.A(count[14]), .B(count[19]), .Z(n29)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i7_2_lut.init = 16'heeee;
    CCU2D add_20292_4 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27753), 
          .COUT(n27754));
    defparam add_20292_4.INIT0 = 16'h5555;
    defparam add_20292_4.INIT1 = 16'h5aaa;
    defparam add_20292_4.INJECT1_0 = "NO";
    defparam add_20292_4.INJECT1_1 = "NO";
    CCU2D add_20292_2 (.A0(count[5]), .B0(count[4]), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27753));
    defparam add_20292_2.INIT0 = 16'h7000;
    defparam add_20292_2.INIT1 = 16'h5aaa;
    defparam add_20292_2.INJECT1_0 = "NO";
    defparam add_20292_2.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27710), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_33.INIT1 = 16'h0000;
    defparam count_2668_add_4_33.INJECT1_0 = "NO";
    defparam count_2668_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27709), .COUT(n27710), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2668_add_4_31.INJECT1_0 = "NO";
    defparam count_2668_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27708), .COUT(n27709), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2668_add_4_29.INJECT1_0 = "NO";
    defparam count_2668_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27707), .COUT(n27708), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2668_add_4_27.INJECT1_0 = "NO";
    defparam count_2668_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27706), .COUT(n27707), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2668_add_4_25.INJECT1_0 = "NO";
    defparam count_2668_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27705), .COUT(n27706), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2668_add_4_23.INJECT1_0 = "NO";
    defparam count_2668_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27704), .COUT(n27705), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2668_add_4_21.INJECT1_0 = "NO";
    defparam count_2668_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27703), .COUT(n27704), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2668_add_4_19.INJECT1_0 = "NO";
    defparam count_2668_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27702), .COUT(n27703), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2668_add_4_17.INJECT1_0 = "NO";
    defparam count_2668_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27701), .COUT(n27702), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2668_add_4_15.INJECT1_0 = "NO";
    defparam count_2668_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27700), .COUT(n27701), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2668_add_4_13.INJECT1_0 = "NO";
    defparam count_2668_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27699), .COUT(n27700), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2668_add_4_11.INJECT1_0 = "NO";
    defparam count_2668_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27698), .COUT(n27699), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2668_add_4_9.INJECT1_0 = "NO";
    defparam count_2668_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27697), .COUT(n27698), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2668_add_4_7.INJECT1_0 = "NO";
    defparam count_2668_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27696), .COUT(n27697), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2668_add_4_5.INJECT1_0 = "NO";
    defparam count_2668_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27695), .COUT(n27696), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2668_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2668_add_4_3.INJECT1_0 = "NO";
    defparam count_2668_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2668_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27695), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668_add_4_1.INIT0 = 16'hF000;
    defparam count_2668_add_4_1.INIT1 = 16'h0555;
    defparam count_2668_add_4_1.INJECT1_0 = "NO";
    defparam count_2668_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2668__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2907), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i1.GSR = "ENABLED";
    FD1S3IX count_2668__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2907), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i2.GSR = "ENABLED";
    FD1S3IX count_2668__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2907), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i3.GSR = "ENABLED";
    FD1S3IX count_2668__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2907), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i4.GSR = "ENABLED";
    FD1S3IX count_2668__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2907), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i5.GSR = "ENABLED";
    FD1S3IX count_2668__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2907), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i6.GSR = "ENABLED";
    FD1S3IX count_2668__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2907), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i7.GSR = "ENABLED";
    FD1S3IX count_2668__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2907), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i8.GSR = "ENABLED";
    FD1S3IX count_2668__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2907), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i9.GSR = "ENABLED";
    FD1S3IX count_2668__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i10.GSR = "ENABLED";
    FD1S3IX count_2668__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i11.GSR = "ENABLED";
    FD1S3IX count_2668__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i12.GSR = "ENABLED";
    FD1S3IX count_2668__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i13.GSR = "ENABLED";
    FD1S3IX count_2668__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i14.GSR = "ENABLED";
    FD1S3IX count_2668__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i15.GSR = "ENABLED";
    FD1S3IX count_2668__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i16.GSR = "ENABLED";
    FD1S3IX count_2668__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i17.GSR = "ENABLED";
    FD1S3IX count_2668__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i18.GSR = "ENABLED";
    FD1S3IX count_2668__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i19.GSR = "ENABLED";
    FD1S3IX count_2668__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i20.GSR = "ENABLED";
    FD1S3IX count_2668__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i21.GSR = "ENABLED";
    FD1S3IX count_2668__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i22.GSR = "ENABLED";
    FD1S3IX count_2668__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i23.GSR = "ENABLED";
    FD1S3IX count_2668__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i24.GSR = "ENABLED";
    FD1S3IX count_2668__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i25.GSR = "ENABLED";
    FD1S3IX count_2668__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i26.GSR = "ENABLED";
    FD1S3IX count_2668__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i27.GSR = "ENABLED";
    FD1S3IX count_2668__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i28.GSR = "ENABLED";
    FD1S3IX count_2668__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i29.GSR = "ENABLED";
    FD1S3IX count_2668__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i30.GSR = "ENABLED";
    FD1S3IX count_2668__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2907), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2668__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ClockDividerP_SP(factor=120000) 
//

module \ClockDividerP_SP(factor=120000)  (debug_c_0, debug_c_c, n34070, 
            n34065, GND_net) /* synthesis syn_module_defined=1 */ ;
    output debug_c_0;
    input debug_c_c;
    input n34070;
    input n34065;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n32167, n20, n19, n21, n28405;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(86[13:18])
    
    wire n2801;
    wire [31:0]n134;
    
    wire n30452, n30148, n30338, n30146, n30298, n30154, n27598, 
        n27597, n27596, n27595, n27594, n27593, n27592, n27591, 
        n27590, n27589, n27588, n27587, n25, n38, n34, n26, 
        n27586, n36, n30, n27585, n27584, n27583, n32, n22;
    
    LUT4 i23121_4_lut_4_lut (.A(n32167), .B(n20), .C(n19), .D(n21), 
         .Z(n28405)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i23121_4_lut_4_lut.init = 16'h0001;
    FD1S3IX clk_o_13 (.D(n28405), .CK(debug_c_c), .CD(n34070), .Q(debug_c_0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(88[9] 107[6])
    defparam clk_o_13.GSR = "ENABLED";
    FD1S3IX count_2660__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2801), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i0.GSR = "ENABLED";
    LUT4 i23052_2_lut (.A(n30452), .B(n34065), .Z(n2801)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23052_2_lut.init = 16'heeee;
    LUT4 i23050_4_lut (.A(n32167), .B(n30148), .C(n30338), .D(n30146), 
         .Z(n30452)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i23050_4_lut.init = 16'h4000;
    LUT4 i22652_2_lut (.A(count[10]), .B(count[12]), .Z(n30148)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22652_2_lut.init = 16'h8888;
    LUT4 i22835_4_lut (.A(count[3]), .B(n30298), .C(n30154), .D(count[0]), 
         .Z(n30338)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22835_4_lut.init = 16'h8000;
    LUT4 i22650_2_lut (.A(count[2]), .B(count[5]), .Z(n30146)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22650_2_lut.init = 16'h8888;
    LUT4 i22795_4_lut (.A(count[1]), .B(count[16]), .C(count[4]), .D(count[15]), 
         .Z(n30298)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22795_4_lut.init = 16'h8000;
    LUT4 i22658_2_lut (.A(count[7]), .B(count[14]), .Z(n30154)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22658_2_lut.init = 16'h8888;
    CCU2D count_2660_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27598), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_33.INIT1 = 16'h0000;
    defparam count_2660_add_4_33.INJECT1_0 = "NO";
    defparam count_2660_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2660_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27597), .COUT(n27598), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2660_add_4_31.INJECT1_0 = "NO";
    defparam count_2660_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2660_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27596), .COUT(n27597), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2660_add_4_29.INJECT1_0 = "NO";
    defparam count_2660_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2660_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27595), .COUT(n27596), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2660_add_4_27.INJECT1_0 = "NO";
    defparam count_2660_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2660_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27594), .COUT(n27595), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2660_add_4_25.INJECT1_0 = "NO";
    defparam count_2660_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2660_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27593), .COUT(n27594), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2660_add_4_23.INJECT1_0 = "NO";
    defparam count_2660_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2660_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27592), .COUT(n27593), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2660_add_4_21.INJECT1_0 = "NO";
    defparam count_2660_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2660_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27591), .COUT(n27592), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2660_add_4_19.INJECT1_0 = "NO";
    defparam count_2660_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2660_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27590), .COUT(n27591), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2660_add_4_17.INJECT1_0 = "NO";
    defparam count_2660_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2660_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27589), .COUT(n27590), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2660_add_4_15.INJECT1_0 = "NO";
    defparam count_2660_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2660_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27588), .COUT(n27589), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2660_add_4_13.INJECT1_0 = "NO";
    defparam count_2660_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2660_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27587), .COUT(n27588), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2660_add_4_11.INJECT1_0 = "NO";
    defparam count_2660_add_4_11.INJECT1_1 = "NO";
    LUT4 i9_4_lut (.A(count[5]), .B(count[16]), .C(count[12]), .D(count[14]), 
         .Z(n21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut_rep_346 (.A(n25), .B(n38), .C(n34), .D(n26), .Z(n32167)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i19_4_lut_rep_346.init = 16'hfffe;
    LUT4 i7_4_lut (.A(count[7]), .B(count[15]), .C(count[4]), .D(count[10]), 
         .Z(n19)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i8_4_lut (.A(count[1]), .B(count[0]), .C(count[2]), .D(count[3]), 
         .Z(n20)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(count[11]), .B(count[13]), .Z(n25)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i5_2_lut.init = 16'heeee;
    CCU2D count_2660_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27586), .COUT(n27587), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2660_add_4_9.INJECT1_0 = "NO";
    defparam count_2660_add_4_9.INJECT1_1 = "NO";
    LUT4 i18_4_lut (.A(count[6]), .B(n36), .C(n30), .D(count[9]), .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i18_4_lut.init = 16'hfffe;
    CCU2D count_2660_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27585), .COUT(n27586), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2660_add_4_7.INJECT1_0 = "NO";
    defparam count_2660_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2660_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27584), .COUT(n27585), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2660_add_4_5.INJECT1_0 = "NO";
    defparam count_2660_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2660_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27583), .COUT(n27584), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2660_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2660_add_4_3.INJECT1_0 = "NO";
    defparam count_2660_add_4_3.INJECT1_1 = "NO";
    LUT4 i14_4_lut (.A(count[20]), .B(count[31]), .C(count[24]), .D(count[30]), 
         .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i14_4_lut.init = 16'hfffe;
    CCU2D count_2660_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27583), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660_add_4_1.INIT0 = 16'hF000;
    defparam count_2660_add_4_1.INIT1 = 16'h0555;
    defparam count_2660_add_4_1.INJECT1_0 = "NO";
    defparam count_2660_add_4_1.INJECT1_1 = "NO";
    LUT4 i6_2_lut (.A(count[21]), .B(count[17]), .Z(n26)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i16_4_lut (.A(count[26]), .B(n32), .C(n22), .D(count[29]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(count[18]), .B(count[28]), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i12_4_lut (.A(count[25]), .B(count[23]), .C(count[8]), .D(count[27]), 
         .Z(n32)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[19]), .B(count[22]), .Z(n22)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(97[9:19])
    defparam i2_2_lut.init = 16'heeee;
    FD1S3IX count_2660__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2801), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i1.GSR = "ENABLED";
    FD1S3IX count_2660__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2801), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i2.GSR = "ENABLED";
    FD1S3IX count_2660__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2801), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i3.GSR = "ENABLED";
    FD1S3IX count_2660__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2801), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i4.GSR = "ENABLED";
    FD1S3IX count_2660__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2801), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i5.GSR = "ENABLED";
    FD1S3IX count_2660__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2801), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i6.GSR = "ENABLED";
    FD1S3IX count_2660__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2801), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i7.GSR = "ENABLED";
    FD1S3IX count_2660__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2801), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i8.GSR = "ENABLED";
    FD1S3IX count_2660__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2801), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i9.GSR = "ENABLED";
    FD1S3IX count_2660__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i10.GSR = "ENABLED";
    FD1S3IX count_2660__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i11.GSR = "ENABLED";
    FD1S3IX count_2660__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i12.GSR = "ENABLED";
    FD1S3IX count_2660__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i13.GSR = "ENABLED";
    FD1S3IX count_2660__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i14.GSR = "ENABLED";
    FD1S3IX count_2660__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i15.GSR = "ENABLED";
    FD1S3IX count_2660__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i16.GSR = "ENABLED";
    FD1S3IX count_2660__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i17.GSR = "ENABLED";
    FD1S3IX count_2660__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i18.GSR = "ENABLED";
    FD1S3IX count_2660__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i19.GSR = "ENABLED";
    FD1S3IX count_2660__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i20.GSR = "ENABLED";
    FD1S3IX count_2660__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i21.GSR = "ENABLED";
    FD1S3IX count_2660__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i22.GSR = "ENABLED";
    FD1S3IX count_2660__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i23.GSR = "ENABLED";
    FD1S3IX count_2660__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i24.GSR = "ENABLED";
    FD1S3IX count_2660__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i25.GSR = "ENABLED";
    FD1S3IX count_2660__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i26.GSR = "ENABLED";
    FD1S3IX count_2660__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i27.GSR = "ENABLED";
    FD1S3IX count_2660__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i28.GSR = "ENABLED";
    FD1S3IX count_2660__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i29.GSR = "ENABLED";
    FD1S3IX count_2660__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i30.GSR = "ENABLED";
    FD1S3IX count_2660__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2801), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(105[16:25])
    defparam count_2660__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module GlobalControlPeripheral
//

module GlobalControlPeripheral (read_value, debug_c_c, n14419, n9478, 
            n34068, read_size, n302, prev_select, \select[1] , n28365, 
            n13412, n34065, n34066, n34070, n34071, \register_addr[0] , 
            \register_addr[1] , timeout_pause, n32285, \register[0][7] , 
            n32227, signal_light_c, rw, n46, n16516, n30075, n16515, 
            n32158, n32200, xbee_pause_c, GND_net, n34067, \databus[1] , 
            n30270, n34069) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    output n14419;
    input n9478;
    input n34068;
    output [2:0]read_size;
    input n302;
    output prev_select;
    input \select[1] ;
    input n28365;
    input n13412;
    input n34065;
    input n34066;
    input n34070;
    input n34071;
    input \register_addr[0] ;
    input \register_addr[1] ;
    input timeout_pause;
    output n32285;
    input \register[0][7] ;
    output n32227;
    output signal_light_c;
    input rw;
    output n46;
    input n16516;
    input n30075;
    input n16515;
    input n32158;
    input n32200;
    input xbee_pause_c;
    input GND_net;
    input n34067;
    input \databus[1] ;
    input n30270;
    input n34069;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]n5914;
    wire [31:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(24[14:22])
    
    wire n14010;
    wire [31:0]n100;
    
    wire prev_clk_1Hz, clk_1Hz;
    wire [31:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(24[14:22])
    
    wire n179;
    wire [31:0]n99;
    
    wire n32271;
    wire [31:0]n271;
    
    wire force_pause, n31919, n31924, n29819, n29820, n29821, n29826, 
        n29822, n29823, n29824, n29825, n29800, n29801, n29802, 
        n29803, n29804, n29805, n29806, n29807, n29808, n29799, 
        n29809, n29810, n29811, n29812, n29813, n29814, n29815, 
        n29816, n29817, n29818, n31920, n31925, n11895, n27342, 
        n27341, n27340, n27339, n27338, n27337, n27336, n27335, 
        n27334, n28876, n27333, n27332, n27331, n27330, n27329, 
        n27328, n27327;
    
    FD1P3IX read_value__i0 (.D(n5914[0]), .SP(n14419), .CD(n9478), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1P3IX uptime_count__i0 (.D(n100[0]), .SP(n14010), .CD(n34068), .CK(debug_c_c), 
            .Q(\register[2] [0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i0.GSR = "ENABLED";
    FD1P3AX read_size_i0_i0 (.D(n302), .SP(n14419), .CK(debug_c_c), .Q(read_size[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_size_i0_i0.GSR = "ENABLED";
    FD1S3AX prev_clk_1Hz_150 (.D(clk_1Hz), .CK(debug_c_c), .Q(prev_clk_1Hz)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam prev_clk_1Hz_150.GSR = "ENABLED";
    FD1S3AX xbee_pause_latched_151 (.D(n179), .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam xbee_pause_latched_151.GSR = "ENABLED";
    FD1S3AX prev_select_149 (.D(\select[1] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam prev_select_149.GSR = "ENABLED";
    LUT4 i15934_4_lut (.A(\register[2] [3]), .B(n9478), .C(n28365), .D(n13412), 
         .Z(n99[3])) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam i15934_4_lut.init = 16'h0323;
    LUT4 i135_2_lut_rep_450 (.A(prev_clk_1Hz), .B(clk_1Hz), .Z(n32271)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(100[9:32])
    defparam i135_2_lut_rep_450.init = 16'h4444;
    LUT4 i2747_2_lut_3_lut (.A(prev_clk_1Hz), .B(clk_1Hz), .C(n34065), 
         .Z(n14010)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(100[9:32])
    defparam i2747_2_lut_3_lut.init = 16'hf4f4;
    FD1P3IX uptime_count__i31 (.D(n100[31]), .SP(n14010), .CD(n34066), 
            .CK(debug_c_c), .Q(\register[2] [31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i31.GSR = "ENABLED";
    FD1P3IX uptime_count__i30 (.D(n100[30]), .SP(n14010), .CD(n34066), 
            .CK(debug_c_c), .Q(\register[2] [30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i30.GSR = "ENABLED";
    FD1P3IX uptime_count__i29 (.D(n100[29]), .SP(n14010), .CD(n34066), 
            .CK(debug_c_c), .Q(\register[2] [29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i29.GSR = "ENABLED";
    FD1P3IX uptime_count__i28 (.D(n100[28]), .SP(n14010), .CD(n34070), 
            .CK(debug_c_c), .Q(\register[2] [28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i28.GSR = "ENABLED";
    FD1P3IX uptime_count__i27 (.D(n100[27]), .SP(n14010), .CD(n34070), 
            .CK(debug_c_c), .Q(\register[2] [27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i27.GSR = "ENABLED";
    FD1P3IX uptime_count__i26 (.D(n100[26]), .SP(n14010), .CD(n34070), 
            .CK(debug_c_c), .Q(\register[2] [26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i26.GSR = "ENABLED";
    FD1P3IX uptime_count__i25 (.D(n100[25]), .SP(n14010), .CD(n34066), 
            .CK(debug_c_c), .Q(\register[2] [25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i25.GSR = "ENABLED";
    FD1P3IX uptime_count__i24 (.D(n100[24]), .SP(n14010), .CD(n34066), 
            .CK(debug_c_c), .Q(\register[2] [24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i24.GSR = "ENABLED";
    FD1P3IX uptime_count__i23 (.D(n100[23]), .SP(n14010), .CD(n34066), 
            .CK(debug_c_c), .Q(\register[2] [23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i23.GSR = "ENABLED";
    FD1P3IX uptime_count__i22 (.D(n100[22]), .SP(n14010), .CD(n34066), 
            .CK(debug_c_c), .Q(\register[2] [22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i22.GSR = "ENABLED";
    FD1P3IX uptime_count__i21 (.D(n100[21]), .SP(n14010), .CD(n34070), 
            .CK(debug_c_c), .Q(\register[2] [21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i21.GSR = "ENABLED";
    FD1P3IX uptime_count__i20 (.D(n100[20]), .SP(n14010), .CD(n34070), 
            .CK(debug_c_c), .Q(\register[2] [20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i20.GSR = "ENABLED";
    FD1P3IX uptime_count__i19 (.D(n100[19]), .SP(n14010), .CD(n34070), 
            .CK(debug_c_c), .Q(\register[2] [19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i19.GSR = "ENABLED";
    FD1P3IX uptime_count__i18 (.D(n100[18]), .SP(n14010), .CD(n34070), 
            .CK(debug_c_c), .Q(\register[2] [18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i18.GSR = "ENABLED";
    FD1P3IX uptime_count__i17 (.D(n100[17]), .SP(n14010), .CD(n34070), 
            .CK(debug_c_c), .Q(\register[2] [17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i17.GSR = "ENABLED";
    FD1P3IX uptime_count__i16 (.D(n100[16]), .SP(n14010), .CD(n34070), 
            .CK(debug_c_c), .Q(\register[2] [16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i16.GSR = "ENABLED";
    FD1P3IX uptime_count__i15 (.D(n271[15]), .SP(n32271), .CD(n34070), 
            .CK(debug_c_c), .Q(\register[2] [15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i15.GSR = "ENABLED";
    FD1P3IX uptime_count__i14 (.D(n271[14]), .SP(n32271), .CD(n34070), 
            .CK(debug_c_c), .Q(\register[2] [14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i14.GSR = "ENABLED";
    FD1P3IX uptime_count__i13 (.D(n271[13]), .SP(n32271), .CD(n34070), 
            .CK(debug_c_c), .Q(\register[2] [13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i13.GSR = "ENABLED";
    FD1P3IX uptime_count__i12 (.D(n271[12]), .SP(n32271), .CD(n34070), 
            .CK(debug_c_c), .Q(\register[2] [12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i12.GSR = "ENABLED";
    FD1P3IX uptime_count__i11 (.D(n271[11]), .SP(n32271), .CD(n34070), 
            .CK(debug_c_c), .Q(\register[2] [11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i11.GSR = "ENABLED";
    FD1P3IX uptime_count__i10 (.D(n271[10]), .SP(n32271), .CD(n34071), 
            .CK(debug_c_c), .Q(\register[2] [10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i10.GSR = "ENABLED";
    FD1P3IX uptime_count__i9 (.D(n271[9]), .SP(n32271), .CD(n34070), .CK(debug_c_c), 
            .Q(\register[2] [9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i9.GSR = "ENABLED";
    FD1P3IX uptime_count__i8 (.D(n271[8]), .SP(n32271), .CD(n34070), .CK(debug_c_c), 
            .Q(\register[2] [8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i8.GSR = "ENABLED";
    FD1P3IX uptime_count__i7 (.D(n271[7]), .SP(n32271), .CD(n34070), .CK(debug_c_c), 
            .Q(\register[2] [7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i7.GSR = "ENABLED";
    FD1P3IX uptime_count__i6 (.D(n271[6]), .SP(n32271), .CD(n34070), .CK(debug_c_c), 
            .Q(\register[2] [6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i6.GSR = "ENABLED";
    FD1P3IX uptime_count__i5 (.D(n100[5]), .SP(n14010), .CD(n34070), .CK(debug_c_c), 
            .Q(\register[2] [5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i5.GSR = "ENABLED";
    FD1P3IX uptime_count__i4 (.D(n100[4]), .SP(n14010), .CD(n34070), .CK(debug_c_c), 
            .Q(\register[2] [4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i4.GSR = "ENABLED";
    FD1P3IX uptime_count__i3 (.D(n100[3]), .SP(n14010), .CD(n34071), .CK(debug_c_c), 
            .Q(\register[2] [3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i3.GSR = "ENABLED";
    FD1P3IX uptime_count__i2 (.D(n271[2]), .SP(n32271), .CD(n34070), .CK(debug_c_c), 
            .Q(\register[2] [2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i2.GSR = "ENABLED";
    FD1P3IX uptime_count__i1 (.D(n271[1]), .SP(n32271), .CD(n34070), .CK(debug_c_c), 
            .Q(\register[2] [1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam uptime_count__i1.GSR = "ENABLED";
    LUT4 register_addr_0__bdd_4_lut_23638 (.A(\register_addr[0] ), .B(force_pause), 
         .C(\register_addr[1] ), .D(\register[2] [1]), .Z(n31919)) /* synthesis lut_function=(!(A (C)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam register_addr_0__bdd_4_lut_23638.init = 16'h5e0e;
    LUT4 i2_3_lut_rep_464 (.A(timeout_pause), .B(force_pause), .C(\register[0] [2]), 
         .Z(n32285)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(39[24:72])
    defparam i2_3_lut_rep_464.init = 16'hfefe;
    LUT4 register_addr_0__bdd_4_lut (.A(\register_addr[0] ), .B(\register[0] [2]), 
         .C(\register_addr[1] ), .D(\register[2] [2]), .Z(n31924)) /* synthesis lut_function=(!(A (C)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam register_addr_0__bdd_4_lut.init = 16'h5e0e;
    LUT4 i14964_2_lut_rep_406_4_lut (.A(timeout_pause), .B(force_pause), 
         .C(\register[0] [2]), .D(\register[0][7] ), .Z(n32227)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(39[24:72])
    defparam i14964_2_lut_rep_406_4_lut.init = 16'h0100;
    LUT4 i14980_2_lut_4_lut (.A(timeout_pause), .B(force_pause), .C(\register[0] [2]), 
         .D(clk_1Hz), .Z(signal_light_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(39[24:72])
    defparam i14980_2_lut_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(\select[1] ), .B(rw), .Z(n46)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(36[19:32])
    defparam i14_2_lut.init = 16'h8888;
    FD1P3IX read_size_i0_i1 (.D(n30075), .SP(n14419), .CD(n16516), .CK(debug_c_c), 
            .Q(read_size[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_size_i0_i1.GSR = "ENABLED";
    FD1P3IX read_size_i0_i2 (.D(n32158), .SP(n14419), .CD(n16515), .CK(debug_c_c), 
            .Q(read_size[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_size_i0_i2.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [4]), 
         .Z(n29819)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_237 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [5]), 
         .Z(n29820)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_237.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_238 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [6]), 
         .Z(n29821)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_238.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_239 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [7]), 
         .Z(n29826)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_239.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_240 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [8]), 
         .Z(n29822)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_240.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_241 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [9]), 
         .Z(n29823)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_241.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_242 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [10]), 
         .Z(n29824)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_242.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_243 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [11]), 
         .Z(n29825)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_243.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_244 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [12]), 
         .Z(n29800)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_244.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_245 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [13]), 
         .Z(n29801)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_245.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_246 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [14]), 
         .Z(n29802)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_246.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_247 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [15]), 
         .Z(n29803)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_247.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_248 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [16]), 
         .Z(n29804)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_248.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_249 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [17]), 
         .Z(n29805)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_249.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_250 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [18]), 
         .Z(n29806)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_250.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_251 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [19]), 
         .Z(n29807)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_251.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_252 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [20]), 
         .Z(n29808)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_252.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_253 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [21]), 
         .Z(n29799)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_253.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_254 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [22]), 
         .Z(n29809)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_254.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_255 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [23]), 
         .Z(n29810)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_255.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_256 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [24]), 
         .Z(n29811)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_256.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_257 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [25]), 
         .Z(n29812)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_257.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_258 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [26]), 
         .Z(n29813)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_258.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_259 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [27]), 
         .Z(n29814)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_259.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_260 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [28]), 
         .Z(n29815)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_260.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_261 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [29]), 
         .Z(n29816)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_261.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_262 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [30]), 
         .Z(n29817)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_262.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_263 (.A(n9478), .B(n28365), .C(n13412), .D(\register[2] [31]), 
         .Z(n29818)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_263.init = 16'h0400;
    LUT4 n1_bdd_2_lut_23639_4_lut (.A(n28365), .B(n9478), .C(n32200), 
         .D(n31919), .Z(n31920)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam n1_bdd_2_lut_23639_4_lut.init = 16'h0200;
    LUT4 n1_bdd_2_lut_23652_4_lut (.A(n28365), .B(n9478), .C(n32200), 
         .D(n31924), .Z(n31925)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam n1_bdd_2_lut_23652_4_lut.init = 16'h0200;
    LUT4 i953_3_lut (.A(prev_select), .B(n34065), .C(\select[1] ), .Z(n14419)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(59[5] 102[8])
    defparam i953_3_lut.init = 16'h1010;
    LUT4 i14928_4_lut (.A(n32200), .B(n28365), .C(n11895), .D(\register_addr[0] ), 
         .Z(n5914[0])) /* synthesis lut_function=(!(A (B)+!A (B ((D)+!C)))) */ ;
    defparam i14928_4_lut.init = 16'h3373;
    LUT4 i5178_3_lut (.A(n32285), .B(\register[2] [0]), .C(\register_addr[1] ), 
         .Z(n11895)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5178_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i3 (.D(n99[3]), .SP(n14419), .CK(debug_c_c), .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3AX read_value__i2 (.D(n31925), .SP(n14419), .CK(debug_c_c), .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3AX read_value__i1 (.D(n31920), .SP(n14419), .CK(debug_c_c), .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i115_1_lut (.A(xbee_pause_c), .Z(n179)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(52[26:39])
    defparam i115_1_lut.init = 16'h5555;
    CCU2D add_135_33 (.A0(\register[2] [31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27342), .S0(n100[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_33.INIT0 = 16'h5aaa;
    defparam add_135_33.INIT1 = 16'h0000;
    defparam add_135_33.INJECT1_0 = "NO";
    defparam add_135_33.INJECT1_1 = "NO";
    CCU2D add_135_31 (.A0(\register[2] [29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27341), .COUT(n27342), .S0(n100[29]), 
          .S1(n100[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_31.INIT0 = 16'h5aaa;
    defparam add_135_31.INIT1 = 16'h5aaa;
    defparam add_135_31.INJECT1_0 = "NO";
    defparam add_135_31.INJECT1_1 = "NO";
    CCU2D add_135_29 (.A0(\register[2] [27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27340), .COUT(n27341), .S0(n100[27]), 
          .S1(n100[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_29.INIT0 = 16'h5aaa;
    defparam add_135_29.INIT1 = 16'h5aaa;
    defparam add_135_29.INJECT1_0 = "NO";
    defparam add_135_29.INJECT1_1 = "NO";
    CCU2D add_135_27 (.A0(\register[2] [25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27339), .COUT(n27340), .S0(n100[25]), 
          .S1(n100[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_27.INIT0 = 16'h5aaa;
    defparam add_135_27.INIT1 = 16'h5aaa;
    defparam add_135_27.INJECT1_0 = "NO";
    defparam add_135_27.INJECT1_1 = "NO";
    FD1P3AX read_value__i4 (.D(n29819), .SP(n14419), .CK(debug_c_c), .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3AX read_value__i5 (.D(n29820), .SP(n14419), .CK(debug_c_c), .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3AX read_value__i6 (.D(n29821), .SP(n14419), .CK(debug_c_c), .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3AX read_value__i7 (.D(n29826), .SP(n14419), .CK(debug_c_c), .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29822), .SP(n14419), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29823), .SP(n14419), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29824), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29825), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29800), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29801), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29802), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29803), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29804), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29805), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29806), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n29807), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29808), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29799), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29809), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29810), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29811), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n29812), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n29813), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n29814), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i27.GSR = "ENABLED";
    CCU2D add_135_25 (.A0(\register[2] [23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27338), .COUT(n27339), .S0(n100[23]), 
          .S1(n100[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_25.INIT0 = 16'h5aaa;
    defparam add_135_25.INIT1 = 16'h5aaa;
    defparam add_135_25.INJECT1_0 = "NO";
    defparam add_135_25.INJECT1_1 = "NO";
    CCU2D add_135_23 (.A0(\register[2] [21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27337), .COUT(n27338), .S0(n100[21]), 
          .S1(n100[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_23.INIT0 = 16'h5aaa;
    defparam add_135_23.INIT1 = 16'h5aaa;
    defparam add_135_23.INJECT1_0 = "NO";
    defparam add_135_23.INJECT1_1 = "NO";
    CCU2D add_135_21 (.A0(\register[2] [19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27336), .COUT(n27337), .S0(n100[19]), 
          .S1(n100[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_21.INIT0 = 16'h5aaa;
    defparam add_135_21.INIT1 = 16'h5aaa;
    defparam add_135_21.INJECT1_0 = "NO";
    defparam add_135_21.INJECT1_1 = "NO";
    FD1P3AX read_value__i28 (.D(n29815), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n29816), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n29817), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n29818), .SP(n14419), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=514, LSE_RLINE=525 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam read_value__i31.GSR = "ENABLED";
    CCU2D add_135_19 (.A0(\register[2] [17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27335), .COUT(n27336), .S0(n100[17]), 
          .S1(n100[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_19.INIT0 = 16'h5aaa;
    defparam add_135_19.INIT1 = 16'h5aaa;
    defparam add_135_19.INJECT1_0 = "NO";
    defparam add_135_19.INJECT1_1 = "NO";
    CCU2D add_135_17 (.A0(\register[2] [15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27334), .COUT(n27335), .S0(n271[15]), 
          .S1(n100[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_17.INIT0 = 16'h5aaa;
    defparam add_135_17.INIT1 = 16'h5aaa;
    defparam add_135_17.INJECT1_0 = "NO";
    defparam add_135_17.INJECT1_1 = "NO";
    FD1P3IX force_pause_152 (.D(\databus[1] ), .SP(n28876), .CD(n34067), 
            .CK(debug_c_c), .Q(force_pause));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(48[9] 103[6])
    defparam force_pause_152.GSR = "ENABLED";
    CCU2D add_135_15 (.A0(\register[2] [13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27333), .COUT(n27334), .S0(n271[13]), 
          .S1(n271[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_15.INIT0 = 16'h5aaa;
    defparam add_135_15.INIT1 = 16'h5aaa;
    defparam add_135_15.INJECT1_0 = "NO";
    defparam add_135_15.INJECT1_1 = "NO";
    CCU2D add_135_13 (.A0(\register[2] [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27332), .COUT(n27333), .S0(n271[11]), 
          .S1(n271[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_13.INIT0 = 16'h5aaa;
    defparam add_135_13.INIT1 = 16'h5aaa;
    defparam add_135_13.INJECT1_0 = "NO";
    defparam add_135_13.INJECT1_1 = "NO";
    CCU2D add_135_11 (.A0(\register[2] [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27331), .COUT(n27332), .S0(n271[9]), .S1(n271[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_11.INIT0 = 16'h5aaa;
    defparam add_135_11.INIT1 = 16'h5aaa;
    defparam add_135_11.INJECT1_0 = "NO";
    defparam add_135_11.INJECT1_1 = "NO";
    CCU2D add_135_9 (.A0(\register[2] [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27330), .COUT(n27331), .S0(n271[7]), .S1(n271[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_9.INIT0 = 16'h5aaa;
    defparam add_135_9.INIT1 = 16'h5aaa;
    defparam add_135_9.INJECT1_0 = "NO";
    defparam add_135_9.INJECT1_1 = "NO";
    CCU2D add_135_7 (.A0(\register[2] [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27329), .COUT(n27330), .S0(n100[5]), .S1(n271[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_7.INIT0 = 16'h5aaa;
    defparam add_135_7.INIT1 = 16'h5aaa;
    defparam add_135_7.INJECT1_0 = "NO";
    defparam add_135_7.INJECT1_1 = "NO";
    CCU2D add_135_5 (.A0(\register[2] [3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27328), .COUT(n27329), .S0(n100[3]), .S1(n100[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_5.INIT0 = 16'h5aaa;
    defparam add_135_5.INIT1 = 16'h5aaa;
    defparam add_135_5.INJECT1_0 = "NO";
    defparam add_135_5.INJECT1_1 = "NO";
    CCU2D add_135_3 (.A0(\register[2] [1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27327), .COUT(n27328), .S0(n271[1]), .S1(n271[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_3.INIT0 = 16'h5aaa;
    defparam add_135_3.INIT1 = 16'h5aaa;
    defparam add_135_3.INJECT1_0 = "NO";
    defparam add_135_3.INJECT1_1 = "NO";
    CCU2D add_135_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\register[2] [0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27327), .S1(n100[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(101[23:39])
    defparam add_135_1.INIT0 = 16'hF000;
    defparam add_135_1.INIT1 = 16'h5555;
    defparam add_135_1.INJECT1_0 = "NO";
    defparam add_135_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(rw), .B(n34065), .C(n30270), .D(\select[1] ), 
         .Z(n28876)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut.init = 16'hcdcc;
    \ClockDividerP(factor=12000000)  uptime_div (.clk_1Hz(clk_1Hz), .debug_c_c(debug_c_c), 
            .n34069(n34069), .GND_net(GND_net), .n34065(n34065)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(105[28] 107[53])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000000) 
//

module \ClockDividerP(factor=12000000)  (clk_1Hz, debug_c_c, n34069, GND_net, 
            n34065) /* synthesis syn_module_defined=1 */ ;
    output clk_1Hz;
    input debug_c_c;
    input n34069;
    input GND_net;
    input n34065;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n7926, n27630;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n134;
    
    wire n27629, n27628, n27627, n27626, n27625, n27624, n27623, 
        n27622, n27621, n27620, n27619, n27618, n27617, n27616, 
        n27615, n2816, n27792, n27791, n27790, n27789, n27788, 
        n27787, n30449, n27, n27804, n25, n26, n24, n19, n32, 
        n28, n20, n27786, n27785, n27784, n27783, n27782, n27781, 
        n29, n26_adj_152;
    
    FD1S3IX clk_o_14 (.D(n7926), .CK(debug_c_c), .CD(n34069), .Q(clk_1Hz));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D count_2661_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27630), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_33.INIT1 = 16'h0000;
    defparam count_2661_add_4_33.INJECT1_0 = "NO";
    defparam count_2661_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27629), .COUT(n27630), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2661_add_4_31.INJECT1_0 = "NO";
    defparam count_2661_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27628), .COUT(n27629), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2661_add_4_29.INJECT1_0 = "NO";
    defparam count_2661_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27627), .COUT(n27628), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2661_add_4_27.INJECT1_0 = "NO";
    defparam count_2661_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27626), .COUT(n27627), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2661_add_4_25.INJECT1_0 = "NO";
    defparam count_2661_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27625), .COUT(n27626), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2661_add_4_23.INJECT1_0 = "NO";
    defparam count_2661_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27624), .COUT(n27625), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2661_add_4_21.INJECT1_0 = "NO";
    defparam count_2661_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27623), .COUT(n27624), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2661_add_4_19.INJECT1_0 = "NO";
    defparam count_2661_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27622), .COUT(n27623), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2661_add_4_17.INJECT1_0 = "NO";
    defparam count_2661_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27621), .COUT(n27622), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2661_add_4_15.INJECT1_0 = "NO";
    defparam count_2661_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27620), .COUT(n27621), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2661_add_4_13.INJECT1_0 = "NO";
    defparam count_2661_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27619), .COUT(n27620), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2661_add_4_11.INJECT1_0 = "NO";
    defparam count_2661_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27618), .COUT(n27619), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2661_add_4_9.INJECT1_0 = "NO";
    defparam count_2661_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27617), .COUT(n27618), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2661_add_4_7.INJECT1_0 = "NO";
    defparam count_2661_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27616), .COUT(n27617), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2661_add_4_5.INJECT1_0 = "NO";
    defparam count_2661_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27615), .COUT(n27616), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2661_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2661_add_4_3.INJECT1_0 = "NO";
    defparam count_2661_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2661_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27615), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661_add_4_1.INIT0 = 16'hF000;
    defparam count_2661_add_4_1.INIT1 = 16'h0555;
    defparam count_2661_add_4_1.INJECT1_0 = "NO";
    defparam count_2661_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2661__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2816), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i0.GSR = "ENABLED";
    CCU2D add_20290_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27792), 
          .S0(n7926));
    defparam add_20290_cout.INIT0 = 16'h0000;
    defparam add_20290_cout.INIT1 = 16'h0000;
    defparam add_20290_cout.INJECT1_0 = "NO";
    defparam add_20290_cout.INJECT1_1 = "NO";
    CCU2D add_20290_24 (.A0(count[30]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[31]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27791), .COUT(n27792));
    defparam add_20290_24.INIT0 = 16'h5555;
    defparam add_20290_24.INIT1 = 16'h5555;
    defparam add_20290_24.INJECT1_0 = "NO";
    defparam add_20290_24.INJECT1_1 = "NO";
    CCU2D add_20290_22 (.A0(count[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[29]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27790), .COUT(n27791));
    defparam add_20290_22.INIT0 = 16'h5555;
    defparam add_20290_22.INIT1 = 16'h5555;
    defparam add_20290_22.INJECT1_0 = "NO";
    defparam add_20290_22.INJECT1_1 = "NO";
    CCU2D add_20290_20 (.A0(count[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27789), .COUT(n27790));
    defparam add_20290_20.INIT0 = 16'h5555;
    defparam add_20290_20.INIT1 = 16'h5555;
    defparam add_20290_20.INJECT1_0 = "NO";
    defparam add_20290_20.INJECT1_1 = "NO";
    CCU2D add_20290_18 (.A0(count[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27788), .COUT(n27789));
    defparam add_20290_18.INIT0 = 16'h5555;
    defparam add_20290_18.INIT1 = 16'h5555;
    defparam add_20290_18.INJECT1_0 = "NO";
    defparam add_20290_18.INJECT1_1 = "NO";
    CCU2D add_20290_16 (.A0(count[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27787), .COUT(n27788));
    defparam add_20290_16.INIT0 = 16'h5aaa;
    defparam add_20290_16.INIT1 = 16'h5555;
    defparam add_20290_16.INJECT1_0 = "NO";
    defparam add_20290_16.INJECT1_1 = "NO";
    LUT4 i23049_2_lut (.A(n30449), .B(n34065), .Z(n2816)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23049_2_lut.init = 16'heeee;
    LUT4 i23047_4_lut (.A(n27), .B(n27804), .C(n25), .D(n26), .Z(n30449)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i23047_4_lut.init = 16'h0004;
    LUT4 i12_4_lut (.A(count[19]), .B(n24), .C(count[8]), .D(count[14]), 
         .Z(n27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(n19), .B(n32), .C(n28), .D(n20), .Z(n27804)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16_4_lut.init = 16'h8000;
    LUT4 i10_4_lut (.A(count[30]), .B(count[22]), .C(count[13]), .D(count[25]), 
         .Z(n25)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i10_4_lut.init = 16'hfffe;
    CCU2D add_20290_14 (.A0(count[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27786), .COUT(n27787));
    defparam add_20290_14.INIT0 = 16'h5aaa;
    defparam add_20290_14.INIT1 = 16'h5555;
    defparam add_20290_14.INJECT1_0 = "NO";
    defparam add_20290_14.INJECT1_1 = "NO";
    CCU2D add_20290_12 (.A0(count[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27785), .COUT(n27786));
    defparam add_20290_12.INIT0 = 16'h5555;
    defparam add_20290_12.INIT1 = 16'h5aaa;
    defparam add_20290_12.INJECT1_0 = "NO";
    defparam add_20290_12.INJECT1_1 = "NO";
    CCU2D add_20290_10 (.A0(count[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27784), .COUT(n27785));
    defparam add_20290_10.INIT0 = 16'h5aaa;
    defparam add_20290_10.INIT1 = 16'h5aaa;
    defparam add_20290_10.INJECT1_0 = "NO";
    defparam add_20290_10.INJECT1_1 = "NO";
    CCU2D add_20290_8 (.A0(count[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27783), .COUT(n27784));
    defparam add_20290_8.INIT0 = 16'h5555;
    defparam add_20290_8.INIT1 = 16'h5aaa;
    defparam add_20290_8.INJECT1_0 = "NO";
    defparam add_20290_8.INJECT1_1 = "NO";
    CCU2D add_20290_6 (.A0(count[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27782), .COUT(n27783));
    defparam add_20290_6.INIT0 = 16'h5555;
    defparam add_20290_6.INIT1 = 16'h5555;
    defparam add_20290_6.INJECT1_0 = "NO";
    defparam add_20290_6.INJECT1_1 = "NO";
    CCU2D add_20290_4 (.A0(count[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27781), .COUT(n27782));
    defparam add_20290_4.INIT0 = 16'h5aaa;
    defparam add_20290_4.INIT1 = 16'h5aaa;
    defparam add_20290_4.INJECT1_0 = "NO";
    defparam add_20290_4.INJECT1_1 = "NO";
    CCU2D add_20290_2 (.A0(count[8]), .B0(count[7]), .C0(GND_net), .D0(GND_net), 
          .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27781));
    defparam add_20290_2.INIT0 = 16'h7000;
    defparam add_20290_2.INIT1 = 16'h5555;
    defparam add_20290_2.INJECT1_0 = "NO";
    defparam add_20290_2.INJECT1_1 = "NO";
    LUT4 i11_4_lut (.A(count[28]), .B(count[15]), .C(count[31]), .D(count[29]), 
         .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut (.A(count[26]), .B(count[24]), .C(count[10]), .D(count[27]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[18]), .B(count[1]), .Z(n19)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i15_4_lut (.A(n29), .B(count[9]), .C(n26_adj_152), .D(count[0]), 
         .Z(n32)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i15_4_lut.init = 16'h8000;
    LUT4 i11_4_lut_adj_235 (.A(count[3]), .B(count[12]), .C(count[5]), 
         .D(count[17]), .Z(n28)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i11_4_lut_adj_235.init = 16'h8000;
    LUT4 i3_2_lut (.A(count[2]), .B(count[11]), .Z(n20)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_236 (.A(count[20]), .B(count[7]), .C(count[23]), 
         .D(count[21]), .Z(n29)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12_4_lut_adj_236.init = 16'h8000;
    LUT4 i9_3_lut (.A(count[16]), .B(count[4]), .C(count[6]), .Z(n26_adj_152)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i9_3_lut.init = 16'h8080;
    FD1S3IX count_2661__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2816), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i1.GSR = "ENABLED";
    FD1S3IX count_2661__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2816), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i2.GSR = "ENABLED";
    FD1S3IX count_2661__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2816), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i3.GSR = "ENABLED";
    FD1S3IX count_2661__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2816), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i4.GSR = "ENABLED";
    FD1S3IX count_2661__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2816), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i5.GSR = "ENABLED";
    FD1S3IX count_2661__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2816), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i6.GSR = "ENABLED";
    FD1S3IX count_2661__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2816), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i7.GSR = "ENABLED";
    FD1S3IX count_2661__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2816), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i8.GSR = "ENABLED";
    FD1S3IX count_2661__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2816), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i9.GSR = "ENABLED";
    FD1S3IX count_2661__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i10.GSR = "ENABLED";
    FD1S3IX count_2661__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i11.GSR = "ENABLED";
    FD1S3IX count_2661__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i12.GSR = "ENABLED";
    FD1S3IX count_2661__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i13.GSR = "ENABLED";
    FD1S3IX count_2661__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i14.GSR = "ENABLED";
    FD1S3IX count_2661__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i15.GSR = "ENABLED";
    FD1S3IX count_2661__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i16.GSR = "ENABLED";
    FD1S3IX count_2661__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i17.GSR = "ENABLED";
    FD1S3IX count_2661__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i18.GSR = "ENABLED";
    FD1S3IX count_2661__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i19.GSR = "ENABLED";
    FD1S3IX count_2661__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i20.GSR = "ENABLED";
    FD1S3IX count_2661__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i21.GSR = "ENABLED";
    FD1S3IX count_2661__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i22.GSR = "ENABLED";
    FD1S3IX count_2661__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i23.GSR = "ENABLED";
    FD1S3IX count_2661__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i24.GSR = "ENABLED";
    FD1S3IX count_2661__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i25.GSR = "ENABLED";
    FD1S3IX count_2661__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i26.GSR = "ENABLED";
    FD1S3IX count_2661__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i27.GSR = "ENABLED";
    FD1S3IX count_2661__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i28.GSR = "ENABLED";
    FD1S3IX count_2661__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i29.GSR = "ENABLED";
    FD1S3IX count_2661__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i30.GSR = "ENABLED";
    FD1S3IX count_2661__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2816), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2661__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module EncoderPeripheral_U11
//

module EncoderPeripheral_U11 (read_value, debug_c_c, n14271, n32160, 
            \read_size[0] , n302, \quadA_delayed[1] , qreset, n6, 
            \quadB_delayed[1] , n13588, n34065, debug_c_0, prev_select, 
            n32182, n32232, n32235, n32278, n9482, \register_addr[0] , 
            encoder_li_c, encoder_lb_c, encoder_la_c, \read_size[2] , 
            n32158, VCC_net, GND_net) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    input n14271;
    input n32160;
    output \read_size[0] ;
    input n302;
    input \quadA_delayed[1] ;
    output qreset;
    input n6;
    input \quadB_delayed[1] ;
    output n13588;
    input n34065;
    input debug_c_0;
    output prev_select;
    input n32182;
    input n32232;
    input n32235;
    input n32278;
    output n9482;
    input \register_addr[0] ;
    input encoder_li_c;
    input encoder_lb_c;
    input encoder_la_c;
    output \read_size[2] ;
    input n32158;
    input VCC_net;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]n100;
    wire [31:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(58[14:22])
    
    wire n29835, n29838, n29849, n29834, n29837, n29836, n29852, 
        n29851, n29842, n29841, n29832, n29840, n29833, n29839, 
        n29846, n29831, n29845, n29830, n29844, n29829, n29843, 
        n29848, n29854, n29855, n29850, n29847, n29828, n29853;
    wire [2:0]quadA_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    
    wire n6_adj_150;
    wire [2:0]quadB_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    
    wire n14779;
    wire [31:0]n180;
    
    FD1P3IX read_value__i0 (.D(n100[0]), .SP(n14271), .CD(n32160), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1P3IX read_size__i1 (.D(n302), .SP(n14271), .CD(n32160), .CK(debug_c_c), 
            .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_size__i1.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(\quadA_delayed[1] ), .B(qreset), .C(n6), .D(\quadB_delayed[1] ), 
         .Z(n13588)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(62[18:35])
    defparam i1_4_lut.init = 16'hedde;
    LUT4 i1_2_lut (.A(n34065), .B(debug_c_0), .Z(qreset)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(62[18:35])
    defparam i1_2_lut.init = 16'heeee;
    FD1S3AX prev_select_126 (.D(n32182), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam prev_select_126.GSR = "ENABLED";
    LUT4 i2_3_lut_3_lut_4_lut (.A(n32232), .B(n32235), .C(n32278), .D(n34065), 
         .Z(n9482)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(77[9:33])
    defparam i2_3_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i1_2_lut_3_lut (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [4]), 
         .Z(n29835)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_207 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [5]), 
         .Z(n29838)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_207.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_208 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [6]), 
         .Z(n29849)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_208.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_209 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [7]), 
         .Z(n29834)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_209.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_210 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [8]), 
         .Z(n29837)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_210.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_211 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [9]), 
         .Z(n29836)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_211.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_212 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [10]), 
         .Z(n29852)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_212.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_213 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [11]), 
         .Z(n29851)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_213.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_214 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [12]), 
         .Z(n29842)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_214.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_215 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [13]), 
         .Z(n29841)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_215.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_216 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [14]), 
         .Z(n29832)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_216.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_217 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [15]), 
         .Z(n29840)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_217.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_218 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [16]), 
         .Z(n29833)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_218.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_219 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [17]), 
         .Z(n29839)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_219.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_220 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [18]), 
         .Z(n29846)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_220.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_221 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [19]), 
         .Z(n29831)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_221.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_222 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [20]), 
         .Z(n29845)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_222.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_223 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [21]), 
         .Z(n29830)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_223.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_224 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [22]), 
         .Z(n29844)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_224.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_225 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [23]), 
         .Z(n29829)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_225.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_226 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [24]), 
         .Z(n29843)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_226.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_227 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [25]), 
         .Z(n29848)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_227.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_228 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [26]), 
         .Z(n29854)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_228.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_229 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [27]), 
         .Z(n29855)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_229.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_230 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [28]), 
         .Z(n29850)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_230.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_231 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [29]), 
         .Z(n29847)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_231.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_232 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [30]), 
         .Z(n29828)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_232.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_233 (.A(\register_addr[0] ), .B(n32160), .C(\register[1] [31]), 
         .Z(n29853)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam i1_2_lut_3_lut_adj_233.init = 16'h2020;
    LUT4 i15021_2_lut (.A(\register[1] [0]), .B(\register_addr[0] ), .Z(n100[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15021_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_234 (.A(quadA_delayed[1]), .B(qreset), .C(n6_adj_150), 
         .D(quadB_delayed[1]), .Z(n14779)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(62[18:35])
    defparam i1_4_lut_adj_234.init = 16'hedde;
    FD1P3IX read_value__i1 (.D(n180[1]), .SP(n14271), .CD(n32160), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n180[2]), .SP(n14271), .CD(n32160), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n180[3]), .SP(n14271), .CD(n32160), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3AX read_value__i4 (.D(n29835), .SP(n14271), .CK(debug_c_c), .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3AX read_value__i5 (.D(n29838), .SP(n14271), .CK(debug_c_c), .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3AX read_value__i6 (.D(n29849), .SP(n14271), .CK(debug_c_c), .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3AX read_value__i7 (.D(n29834), .SP(n14271), .CK(debug_c_c), .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29837), .SP(n14271), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29836), .SP(n14271), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29852), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29851), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29842), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29841), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29832), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29840), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29833), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29839), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29846), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n29831), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29845), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29830), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29844), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29829), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29843), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n29848), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n29854), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n29855), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n29850), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n29847), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n29828), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n29853), .SP(n14271), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i31.GSR = "ENABLED";
    LUT4 mux_115_Mux_1_i1_3_lut (.A(encoder_li_c), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n180[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_2_i1_3_lut (.A(encoder_lb_c), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n180[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_3_i1_3_lut (.A(encoder_la_c), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n180[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_3_i1_3_lut.init = 16'hcaca;
    FD1P3IX read_size__i2 (.D(n32158), .SP(n14271), .CD(n32160), .CK(debug_c_c), 
            .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=671, LSE_RLINE=681 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_size__i2.GSR = "ENABLED";
    QuadratureDecoder_U6 q (.\register[1] ({\register[1] }), .debug_c_c(debug_c_c), 
            .qreset(qreset), .VCC_net(VCC_net), .GND_net(GND_net), .encoder_lb_c(encoder_lb_c), 
            .n14779(n14779), .encoder_la_c(encoder_la_c), .\quadB_delayed[1] (quadB_delayed[1]), 
            .\quadA_delayed[1] (quadA_delayed[1]), .n6(n6_adj_150)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(92[20] 96[37])
    
endmodule
//
// Verilog Description of module QuadratureDecoder_U6
//

module QuadratureDecoder_U6 (\register[1] , debug_c_c, qreset, VCC_net, 
            GND_net, encoder_lb_c, n14779, encoder_la_c, \quadB_delayed[1] , 
            \quadA_delayed[1] , n6) /* synthesis syn_module_defined=1 */ ;
    output [31:0]\register[1] ;
    input debug_c_c;
    input qreset;
    input VCC_net;
    input GND_net;
    input encoder_lb_c;
    input n14779;
    input encoder_la_c;
    output \quadB_delayed[1] ;
    output \quadA_delayed[1] ;
    output n6;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(15[13:18])
    wire [2:0]quadB_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    wire [31:0]n100;
    wire [2:0]quadA_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    wire [31:0]n4298;
    
    wire n27065, n27064, n27063, n27062, n27061, n27060, n27059, 
        n27058, n27057, n27056, n27050, n27055, n27054, n27053, 
        n27052, n27051;
    
    FD1P3AX count_at_reset_i0_i0 (.D(count[0]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i0.GSR = "ENABLED";
    IFS1P3DX quadB_delayed_i0 (.D(encoder_lb_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadB_delayed[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i0.GSR = "ENABLED";
    FD1P3IX count__i0 (.D(n100[0]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i0.GSR = "ENABLED";
    IFS1P3DX quadA_delayed_i0 (.D(encoder_la_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadA_delayed[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i0.GSR = "ENABLED";
    FD1P3IX count__i31 (.D(n4298[31]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i31.GSR = "ENABLED";
    FD1P3IX count__i30 (.D(n4298[30]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i30.GSR = "ENABLED";
    FD1P3IX count__i29 (.D(n4298[29]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i29.GSR = "ENABLED";
    FD1P3IX count__i28 (.D(n4298[28]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i28.GSR = "ENABLED";
    FD1P3IX count__i27 (.D(n4298[27]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i27.GSR = "ENABLED";
    FD1P3IX count__i26 (.D(n4298[26]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i26.GSR = "ENABLED";
    FD1P3IX count__i25 (.D(n4298[25]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i25.GSR = "ENABLED";
    FD1P3IX count__i24 (.D(n4298[24]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i24.GSR = "ENABLED";
    FD1P3IX count__i23 (.D(n4298[23]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i23.GSR = "ENABLED";
    FD1P3IX count__i22 (.D(n4298[22]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i22.GSR = "ENABLED";
    FD1P3IX count__i21 (.D(n4298[21]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i21.GSR = "ENABLED";
    FD1P3IX count__i20 (.D(n4298[20]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i20.GSR = "ENABLED";
    FD1P3IX count__i19 (.D(n4298[19]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i19.GSR = "ENABLED";
    FD1P3IX count__i18 (.D(n4298[18]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i18.GSR = "ENABLED";
    FD1P3IX count__i17 (.D(n4298[17]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i17.GSR = "ENABLED";
    FD1P3IX count__i16 (.D(n4298[16]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i16.GSR = "ENABLED";
    FD1P3IX count__i15 (.D(n4298[15]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i15.GSR = "ENABLED";
    FD1P3IX count__i14 (.D(n4298[14]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i14.GSR = "ENABLED";
    FD1P3IX count__i13 (.D(n4298[13]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i13.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n4298[12]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i12.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n4298[11]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n4298[10]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n4298[9]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n4298[8]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n4298[7]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n4298[6]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n4298[5]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n4298[4]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n4298[3]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n4298[2]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n4298[1]), .SP(n14779), .CD(qreset), .CK(debug_c_c), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i1.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i1 (.D(count[1]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i1.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i2 (.D(count[2]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i2.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i3 (.D(count[3]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i3.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i4 (.D(count[4]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i4.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i5 (.D(count[5]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i5.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i6 (.D(count[6]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i6.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i7 (.D(count[7]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i7.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i8 (.D(count[8]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i8.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i9 (.D(count[9]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i9.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i10 (.D(count[10]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i10.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i11 (.D(count[11]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i11.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i12 (.D(count[12]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i12.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i13 (.D(count[13]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i13.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i14 (.D(count[14]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i14.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i15 (.D(count[15]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i15.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i16 (.D(count[16]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i16.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i17 (.D(count[17]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i17.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i18 (.D(count[18]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i18.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i19 (.D(count[19]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i19.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i20 (.D(count[20]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i20.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i21 (.D(count[21]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i21.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i22 (.D(count[22]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i22.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i23 (.D(count[23]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i23.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i24 (.D(count[24]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i24.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i25 (.D(count[25]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i25.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i26 (.D(count[26]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i26.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i27 (.D(count[27]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i27.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i28 (.D(count[28]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i28.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i29 (.D(count[29]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i29.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i30 (.D(count[30]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i30.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i31 (.D(count[31]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i31.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i1 (.D(quadB_delayed[0]), .CK(debug_c_c), .Q(\quadB_delayed[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i1.GSR = "ENABLED";
    CCU2D add_1672_33 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[30]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[31]), .D1(GND_net), .CIN(n27065), .S0(n4298[30]), 
          .S1(n4298[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_33.INIT0 = 16'h6969;
    defparam add_1672_33.INIT1 = 16'h6969;
    defparam add_1672_33.INJECT1_0 = "NO";
    defparam add_1672_33.INJECT1_1 = "NO";
    FD1S3AX quadB_delayed_i2 (.D(\quadB_delayed[1] ), .CK(debug_c_c), .Q(quadB_delayed[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i2.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i1 (.D(quadA_delayed[0]), .CK(debug_c_c), .Q(\quadA_delayed[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i2 (.D(\quadA_delayed[1] ), .CK(debug_c_c), .Q(quadA_delayed[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i2.GSR = "ENABLED";
    CCU2D add_1672_31 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[28]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[29]), .D1(GND_net), .CIN(n27064), .COUT(n27065), 
          .S0(n4298[28]), .S1(n4298[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_31.INIT0 = 16'h6969;
    defparam add_1672_31.INIT1 = 16'h6969;
    defparam add_1672_31.INJECT1_0 = "NO";
    defparam add_1672_31.INJECT1_1 = "NO";
    CCU2D add_1672_29 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[26]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[27]), .D1(GND_net), .CIN(n27063), .COUT(n27064), 
          .S0(n4298[26]), .S1(n4298[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_29.INIT0 = 16'h6969;
    defparam add_1672_29.INIT1 = 16'h6969;
    defparam add_1672_29.INJECT1_0 = "NO";
    defparam add_1672_29.INJECT1_1 = "NO";
    CCU2D add_1672_27 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[24]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[25]), .D1(GND_net), .CIN(n27062), .COUT(n27063), 
          .S0(n4298[24]), .S1(n4298[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_27.INIT0 = 16'h6969;
    defparam add_1672_27.INIT1 = 16'h6969;
    defparam add_1672_27.INJECT1_0 = "NO";
    defparam add_1672_27.INJECT1_1 = "NO";
    CCU2D add_1672_25 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[22]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[23]), .D1(GND_net), .CIN(n27061), .COUT(n27062), 
          .S0(n4298[22]), .S1(n4298[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_25.INIT0 = 16'h6969;
    defparam add_1672_25.INIT1 = 16'h6969;
    defparam add_1672_25.INJECT1_0 = "NO";
    defparam add_1672_25.INJECT1_1 = "NO";
    CCU2D add_1672_23 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[20]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[21]), .D1(GND_net), .CIN(n27060), .COUT(n27061), 
          .S0(n4298[20]), .S1(n4298[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_23.INIT0 = 16'h6969;
    defparam add_1672_23.INIT1 = 16'h6969;
    defparam add_1672_23.INJECT1_0 = "NO";
    defparam add_1672_23.INJECT1_1 = "NO";
    CCU2D add_1672_21 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[18]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[19]), .D1(GND_net), .CIN(n27059), .COUT(n27060), 
          .S0(n4298[18]), .S1(n4298[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_21.INIT0 = 16'h6969;
    defparam add_1672_21.INIT1 = 16'h6969;
    defparam add_1672_21.INJECT1_0 = "NO";
    defparam add_1672_21.INJECT1_1 = "NO";
    CCU2D add_1672_19 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[16]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[17]), .D1(GND_net), .CIN(n27058), .COUT(n27059), 
          .S0(n4298[16]), .S1(n4298[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_19.INIT0 = 16'h6969;
    defparam add_1672_19.INIT1 = 16'h6969;
    defparam add_1672_19.INJECT1_0 = "NO";
    defparam add_1672_19.INJECT1_1 = "NO";
    CCU2D add_1672_17 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[14]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[15]), .D1(GND_net), .CIN(n27057), .COUT(n27058), 
          .S0(n4298[14]), .S1(n4298[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_17.INIT0 = 16'h6969;
    defparam add_1672_17.INIT1 = 16'h6969;
    defparam add_1672_17.INJECT1_0 = "NO";
    defparam add_1672_17.INJECT1_1 = "NO";
    CCU2D add_1672_15 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[12]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[13]), .D1(GND_net), .CIN(n27056), .COUT(n27057), 
          .S0(n4298[12]), .S1(n4298[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_15.INIT0 = 16'h6969;
    defparam add_1672_15.INIT1 = 16'h6969;
    defparam add_1672_15.INJECT1_0 = "NO";
    defparam add_1672_15.INJECT1_1 = "NO";
    CCU2D add_1672_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27050));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_1.INIT0 = 16'hF000;
    defparam add_1672_1.INIT1 = 16'h6666;
    defparam add_1672_1.INJECT1_0 = "NO";
    defparam add_1672_1.INJECT1_1 = "NO";
    CCU2D add_1672_13 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[10]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[11]), .D1(GND_net), .CIN(n27055), .COUT(n27056), 
          .S0(n4298[10]), .S1(n4298[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_13.INIT0 = 16'h6969;
    defparam add_1672_13.INIT1 = 16'h6969;
    defparam add_1672_13.INJECT1_0 = "NO";
    defparam add_1672_13.INJECT1_1 = "NO";
    CCU2D add_1672_11 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[8]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[9]), .D1(GND_net), .CIN(n27054), .COUT(n27055), 
          .S0(n4298[8]), .S1(n4298[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_11.INIT0 = 16'h6969;
    defparam add_1672_11.INIT1 = 16'h6969;
    defparam add_1672_11.INJECT1_0 = "NO";
    defparam add_1672_11.INJECT1_1 = "NO";
    LUT4 i2_2_lut (.A(quadB_delayed[2]), .B(quadA_delayed[2]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(18[22:95])
    defparam i2_2_lut.init = 16'h6666;
    CCU2D add_1672_9 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[6]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[7]), .D1(GND_net), .CIN(n27053), .COUT(n27054), 
          .S0(n4298[6]), .S1(n4298[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_9.INIT0 = 16'h6969;
    defparam add_1672_9.INIT1 = 16'h6969;
    defparam add_1672_9.INJECT1_0 = "NO";
    defparam add_1672_9.INJECT1_1 = "NO";
    CCU2D add_1672_7 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[4]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[5]), .D1(GND_net), .CIN(n27052), .COUT(n27053), 
          .S0(n4298[4]), .S1(n4298[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_7.INIT0 = 16'h6969;
    defparam add_1672_7.INIT1 = 16'h6969;
    defparam add_1672_7.INJECT1_0 = "NO";
    defparam add_1672_7.INJECT1_1 = "NO";
    CCU2D add_1672_5 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[2]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[3]), .D1(GND_net), .CIN(n27051), .COUT(n27052), 
          .S0(n4298[2]), .S1(n4298[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_5.INIT0 = 16'h6969;
    defparam add_1672_5.INIT1 = 16'h6969;
    defparam add_1672_5.INJECT1_0 = "NO";
    defparam add_1672_5.INJECT1_1 = "NO";
    CCU2D add_1672_3 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[0]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[1]), .D1(GND_net), .CIN(n27050), .COUT(n27051), 
          .S0(n100[0]), .S1(n4298[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1672_3.INIT0 = 16'h9696;
    defparam add_1672_3.INIT1 = 16'h6969;
    defparam add_1672_3.INJECT1_0 = "NO";
    defparam add_1672_3.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \ProtocolInterface(baud_div=12) 
//

module \ProtocolInterface(baud_div=12)  (register_addr, debug_c_c, n13118, 
            n29983, databus, n224, n3862, debug_c_7, n32213, n32261, 
            n32235, n32315, n29712, \select[5] , rw, n19559, n32152, 
            n34064, n13567, databus_out, \sendcount[1] , n32153, n224_adj_56, 
            n3948, n32172, n32278, n34065, n13560, \select[7] , 
            \select[4] , \select[3] , \select[2] , \select[1] , n1432, 
            n13545, prev_select, n2760, n32279, n29750, n32154, 
            n13885, n21718, n32282, n32233, n32202, n32231, n32137, 
            n32253, n112, n30075, debug_c_5, n32251, n52, prev_select_adj_41, 
            n32181, n32305, n32182, n29713, n32178, n5774, n32314, 
            n28302, n32316, n32252, n13576, n13899, n32165, n13769, 
            \control_reg[7] , n8585, n32168, prev_select_adj_42, n32163, 
            n32140, n29977, n4034, n64, \control_reg[7]_adj_43 , n8594, 
            \control_reg[7]_adj_44 , n1, n12746, n13, n18, n14, 
            n32155, \reg_size[2] , n32284, n28062, n32285, n34, 
            n28053, n32, debug_c_2, debug_c_3, debug_c_4, \steps_reg[5] , 
            n14_adj_45, n28049, \control_reg[7]_adj_46 , n32_adj_47, 
            \steps_reg[6] , n13_adj_48, \steps_reg[3] , n12, n4, n28061, 
            n32_adj_49, \steps_reg[5]_adj_50 , n14_adj_51, \steps_reg[6]_adj_52 , 
            n13_adj_53, n32234, n13412, \steps_reg[3]_adj_54 , n12_adj_55, 
            n8576, \reset_count[14] , \reset_count[13] , \reset_count[12] , 
            n29954, uart_tx_c, GND_net, uart_rx_c) /* synthesis syn_module_defined=1 */ ;
    output [7:0]register_addr;
    input debug_c_c;
    input n13118;
    output n29983;
    input [31:0]databus;
    input [31:0]n224;
    output [31:0]n3862;
    output debug_c_7;
    output n32213;
    output n32261;
    output n32235;
    input n32315;
    output n29712;
    output \select[5] ;
    output rw;
    output n19559;
    input n32152;
    output n34064;
    input n13567;
    output [31:0]databus_out;
    output \sendcount[1] ;
    input n32153;
    input [31:0]n224_adj_56;
    output [31:0]n3948;
    input n32172;
    output n32278;
    input n34065;
    output n13560;
    output \select[7] ;
    output \select[4] ;
    output \select[3] ;
    output \select[2] ;
    output \select[1] ;
    output n1432;
    output n13545;
    input prev_select;
    output n2760;
    output n32279;
    input n29750;
    input n32154;
    output n13885;
    output n21718;
    output n32282;
    output n32233;
    output n32202;
    output n32231;
    output n32137;
    input n32253;
    output n112;
    output n30075;
    output debug_c_5;
    input n32251;
    output n52;
    input prev_select_adj_41;
    output n32181;
    output n32305;
    output n32182;
    output n29713;
    output n32178;
    output n5774;
    output n32314;
    output n28302;
    output n32316;
    output n32252;
    input n13576;
    output n13899;
    input n32165;
    output n13769;
    input \control_reg[7] ;
    output n8585;
    output n32168;
    input prev_select_adj_42;
    output n32163;
    output n32140;
    input n29977;
    output n4034;
    output n64;
    input \control_reg[7]_adj_43 ;
    output n8594;
    input \control_reg[7]_adj_44 ;
    output n1;
    input n12746;
    input n13;
    input n18;
    input n14;
    output n32155;
    input \reg_size[2] ;
    input n32284;
    input n28062;
    input n32285;
    output n34;
    input n28053;
    output n32;
    output debug_c_2;
    output debug_c_3;
    output debug_c_4;
    input \steps_reg[5] ;
    output n14_adj_45;
    input n28049;
    input \control_reg[7]_adj_46 ;
    output n32_adj_47;
    input \steps_reg[6] ;
    output n13_adj_48;
    input \steps_reg[3] ;
    output n12;
    output n4;
    input n28061;
    output n32_adj_49;
    input \steps_reg[5]_adj_50 ;
    output n14_adj_51;
    input \steps_reg[6]_adj_52 ;
    output n13_adj_53;
    input n32234;
    output n13412;
    input \steps_reg[3]_adj_54 ;
    output n12_adj_55;
    output n8576;
    input \reset_count[14] ;
    input \reset_count[13] ;
    input \reset_count[12] ;
    input n29954;
    output uart_tx_c;
    input GND_net;
    input uart_rx_c;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(455[15:21])
    
    wire n2746;
    wire [7:0]\buffer[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire escape, n12924, n6;
    wire [31:0]n1414;
    
    wire n10915;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(52[12:19])
    
    wire n32180, n16522;
    wire [7:0]esc_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(51[12:20])
    
    wire n29552;
    wire [7:0]rx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(50[13:20])
    
    wire n13_c;
    wire [7:0]\buffer[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n30012, n16289, n1867, n32122;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    
    wire n32177, n32156, n22501, n15653;
    wire [3:0]n1810;
    
    wire n1815, n15654, n15626, n32123;
    wire [7:0]n2156;
    wire [3:0]bufcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(46[12:20])
    
    wire n32169, n15360, n31123, n2748;
    wire [7:0]\buffer[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n9;
    wire [4:0]n9281;
    
    wire n15359, n28238, n10136, n30294, n30083, n15661, n32120, 
        n16363, n32121, n13422, n21572, n34073, n29226, n32268, 
        n32223, n32269;
    wire [7:0]\buffer[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]\buffer[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n31121, n32_c, n32322, n32326;
    wire [7:0]\buffer[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n32325, n32329, n32328, n15625, n15641, n16519;
    wire [7:0]n9241;
    
    wire n32275, n32332, n32331, n32229;
    wire [7:0]n5765;
    
    wire n32321, n34061, n32335, n32334, n32276, n32338, n32337, 
        n32341, n32340, n32344, n32343, n32347, n32346, n29532, 
        n9_adj_38, n32397, n29702, n32280, n32395, n14_c, n29720, 
        n29727, n29721, n29725, n29723, n29719, n29728, n29726, 
        n29724, n29722, n29731, n29729, n29735, n29732, n29715, 
        n29730, n32201, n29733, n32281, n29716, n32230, n7, n29739, 
        n29737, n29736, n14_adj_39, n29734, n29742, n29741, n29738, 
        n29745, n29740, n29743, n29744, n29717, n29746, n29718, 
        send, n28225, n12484, n32289, n31812, n31813, n30052, 
        n30053, n32291, n15624, n28639, n32239, n30023, n30022, 
        n32292, n31814, n31815, n29547, n28299, n32333, n31122, 
        n4_c, n32345, n4_adj_44, n32342, n4_adj_45, n32336, n4_adj_46, 
        n32348, n4_adj_47, n32327, n4_adj_48, n32330, n13115, n1519, 
        n4_adj_49, n32339, n15640, n10, n8, n29368, n15, n29707, 
        n6_adj_52, n13034, n29645, n29276, n30328, n11, n11_adj_54, 
        n11_adj_55, n11_adj_56, n11_adj_57, n11928, n29575, n29634, 
        n30284, n31805, n11_adj_58, n11_adj_59, n11_adj_60, n11_adj_61, 
        n11_adj_62, n11_adj_63, n11_adj_64, n11_adj_65, n11_adj_66, 
        n11_adj_67, n11_adj_68, busy, n1525, n1526, n2687, n11158, 
        n11930, n29924, n31117, n35, n29278, n11151, n11932, n29244, 
        n29204, n29202, n32319, n32320, n29218, n29208, n5, n28156, 
        n29903, n29200, n29214, n29210, n29224, n29242, n29216, 
        n29220, n29222, n29228, n29230, n30316, n9411, n5_adj_73, 
        n28134, n5_adj_74, n28136, n5_adj_75, n28104, n5_adj_76, 
        n28106, n5_adj_77, n28137, n5_adj_78, n28143, n5_adj_79, 
        n28147, n5_adj_80, n28145, n5_adj_81, n28146, n5_adj_82, 
        n28142, n5_adj_83, n28149, n5_adj_84, n28153, n5_adj_85, 
        n28150, n5_adj_86, n28152, n5_adj_87, n28151, n5_adj_88, 
        n28148, n5_adj_89, n28154, n5_adj_91, n28157, n5_adj_92, 
        n28161, n5_adj_93, n28105, n5_adj_94, n28172, n5_adj_95, 
        n28162, n5_adj_96, n28168, n5_adj_97, n28163, n5_adj_98, 
        n28169, n5_adj_100, n28165, n5_adj_101, n28171, n5_adj_103, 
        n28166, n5_adj_104, n28170, n5_adj_105, n28167, n5_adj_106, 
        n28160, n7_adj_107, n1_adj_113, n6_adj_114, n29701, n27934, 
        n32323, n8_adj_125, n8_adj_126, n6_adj_127;
    wire [3:0]n9547;
    
    FD1P3AX reg_addr_i0_i0 (.D(\buffer[1] [0]), .SP(n2746), .CK(debug_c_c), 
            .Q(register_addr[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i0.GSR = "ENABLED";
    LUT4 mux_1542_i27_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[26]), 
         .D(n224[26]), .Z(n3862[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i27_3_lut_4_lut.init = 16'hf780;
    LUT4 i9017_4_lut (.A(escape), .B(n12924), .C(n6), .D(n1414[3]), 
         .Z(n10915)) /* synthesis lut_function=(!(A (C (D))+!A (B+!(C (D))))) */ ;
    defparam i9017_4_lut.init = 16'h1aaa;
    LUT4 i2_2_lut (.A(debug_c_7), .B(n32213), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    FD1P3IX tx_data_i0_i2 (.D(esc_data[2]), .SP(n32180), .CD(n16522), 
            .CK(debug_c_c), .Q(tx_data[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_440 (.A(register_addr[5]), .B(register_addr[4]), .Z(n32261)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_440.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(register_addr[4]), 
         .C(n32235), .D(n32315), .Z(n29712)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0008;
    FD1P3IX tx_data_i0_i5 (.D(esc_data[5]), .SP(n32180), .CD(n16522), 
            .CK(debug_c_c), .Q(tx_data[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(\select[5] ), .B(rw), .Z(n19559)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(register_addr[4]), .B(n32152), .C(register_addr[5]), 
         .D(n34064), .Z(n29983)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_4_lut.init = 16'h0080;
    LUT4 i2_4_lut (.A(n29552), .B(rx_data[4]), .C(rx_data[1]), .D(rx_data[3]), 
         .Z(n12924)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'hbfff;
    LUT4 i2_4_lut_adj_51 (.A(n13_c), .B(rx_data[5]), .C(rx_data[2]), .D(rx_data[0]), 
         .Z(n29552)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i2_4_lut_adj_51.init = 16'hfeff;
    LUT4 equal_142_i13_2_lut (.A(rx_data[6]), .B(rx_data[7]), .Z(n13_c)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(134[12:17])
    defparam equal_142_i13_2_lut.init = 16'heeee;
    LUT4 mux_1542_i26_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[25]), 
         .D(n224[25]), .Z(n3862[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i26_3_lut_4_lut.init = 16'hf780;
    LUT4 \buffer_0[[0__bdd_4_lut_23736  (.A(\buffer[0] [0]), .B(n30012), 
         .C(n16289), .D(n1867), .Z(n32122)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;
    defparam \buffer_0[[0__bdd_4_lut_23736 .init = 16'h11f0;
    FD1P3IX sendcount__i0 (.D(n22501), .SP(n32177), .CD(n32156), .CK(debug_c_c), 
            .Q(sendcount[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i0.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i6 (.D(esc_data[6]), .SP(n32180), .CD(n16522), 
            .CK(debug_c_c), .Q(tx_data[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    LUT4 mux_1542_i25_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[24]), 
         .D(n224[24]), .Z(n3862[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i25_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1542_i24_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[23]), 
         .D(n224[23]), .Z(n3862[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i24_3_lut_4_lut.init = 16'hf780;
    PFUMX i8933 (.BLUT(n15653), .ALUT(n1810[1]), .C0(n1815), .Z(n15654));
    LUT4 mux_1542_i23_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[22]), 
         .D(n224[22]), .Z(n3862[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 \buffer_0[[0__bdd_4_lut  (.A(\buffer[0] [0]), .B(n30012), .C(n15626), 
         .D(n1867), .Z(n32123)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C))) */ ;
    defparam \buffer_0[[0__bdd_4_lut .init = 16'h22f0;
    FD1P3AX tx_data_i0_i0 (.D(n2156[0]), .SP(n32180), .CK(debug_c_c), 
            .Q(tx_data[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    FD1S3IX bufcount__i0 (.D(n15360), .CK(debug_c_c), .CD(n32169), .Q(bufcount[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i0.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i0 (.D(n31123), .SP(n13567), .CK(debug_c_c), .Q(esc_data[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i0.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i0 (.D(\buffer[2] [0]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i0.GSR = "ENABLED";
    LUT4 i15125_3_lut_4_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(n9), 
         .D(sendcount[2]), .Z(n9281[2])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C))) */ ;
    defparam i15125_3_lut_4_lut.init = 16'h7f8f;
    PFUMX i8639 (.BLUT(n15359), .ALUT(n28238), .C0(n1815), .Z(n15360));
    LUT4 i3394_2_lut_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(sendcount[2]), 
         .Z(n10136)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i3394_2_lut_3_lut.init = 16'h8080;
    LUT4 i22791_3_lut_4_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(sendcount[3]), 
         .D(sendcount[2]), .Z(n30294)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22791_3_lut_4_lut.init = 16'h8000;
    LUT4 \buffer_0[[1__bdd_4_lut_23735  (.A(\buffer[0] [1]), .B(n30083), 
         .C(n15661), .D(n1867), .Z(n32120)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;
    defparam \buffer_0[[1__bdd_4_lut_23735 .init = 16'h11f0;
    LUT4 \buffer_0[[1__bdd_4_lut  (.A(\buffer[0] [1]), .B(n30083), .C(n16363), 
         .D(n1867), .Z(n32121)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C))) */ ;
    defparam \buffer_0[[1__bdd_4_lut .init = 16'h22f0;
    FD1S3JX state_FSM_i1 (.D(n13422), .CK(debug_c_c), .PD(n32169), .Q(n1414[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i1.GSR = "ENABLED";
    FD1P3IX buffer_0___i1 (.D(n29226), .SP(n21572), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[0] [0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i1.GSR = "ENABLED";
    LUT4 mux_1542_i22_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[21]), 
         .D(n224[21]), .Z(n3862[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1542_i21_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[20]), 
         .D(n224[20]), .Z(n3862[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 i14936_2_lut_rep_447 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n32268)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14936_2_lut_rep_447.init = 16'heeee;
    LUT4 mux_1542_i20_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[19]), 
         .D(n224[19]), .Z(n3862[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1542_i19_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[18]), 
         .D(n224[18]), .Z(n3862[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_402_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(sendcount[2]), 
         .Z(n32223)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam i1_2_lut_rep_402_3_lut.init = 16'h1e1e;
    LUT4 i3385_2_lut_rep_448 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n32269)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i3385_2_lut_rep_448.init = 16'h9999;
    LUT4 n12742_bdd_4_lut_23350_4_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(\buffer[5] [0]), .D(\buffer[4] [0]), .Z(n31121)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam n12742_bdd_4_lut_23350_4_lut.init = 16'h6420;
    LUT4 i15126_2_lut_2_lut_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(n9), .Z(n9281[1])) /* synthesis lut_function=(!(A (B (C))+!A !(B+!(C)))) */ ;
    defparam i15126_2_lut_2_lut_3_lut.init = 16'h6f6f;
    LUT4 mux_1564_i20_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[19]), 
         .D(n224_adj_56[19]), .Z(n3948[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 i42_4_lut_4_lut (.A(esc_data[4]), .B(esc_data[1]), .C(esc_data[3]), 
         .D(esc_data[2]), .Z(n32_c)) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A (B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i42_4_lut_4_lut.init = 16'h0881;
    LUT4 i1_4_lut_else_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(\sendcount[1] ), 
         .D(sendcount[2]), .Z(n32322)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h4001;
    LUT4 mux_1564_i19_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[18]), 
         .D(n224_adj_56[18]), .Z(n3948[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_52 (.A(n32172), .B(n32278), .C(n34065), 
         .D(register_addr[0]), .Z(n13560)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_52.init = 16'hf0f4;
    LUT4 i22877_then_3_lut (.A(\buffer[0] [6]), .B(\buffer[2] [6]), .C(\sendcount[1] ), 
         .Z(n32326)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22877_then_3_lut.init = 16'hcaca;
    LUT4 i22877_else_3_lut (.A(\buffer[3] [6]), .B(\buffer[1] [6]), .C(\sendcount[1] ), 
         .Z(n32325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22877_else_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i18_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[17]), 
         .D(n224_adj_56[17]), .Z(n3948[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i18_3_lut_4_lut.init = 16'hf780;
    FD1P3IX tx_data_i0_i7 (.D(esc_data[7]), .SP(n32180), .CD(n16522), 
            .CK(debug_c_c), .Q(tx_data[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    LUT4 i22880_then_3_lut (.A(\buffer[0] [5]), .B(\buffer[2] [5]), .C(\sendcount[1] ), 
         .Z(n32329)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22880_then_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i17_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[16]), 
         .D(n224_adj_56[16]), .Z(n3948[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i22880_else_3_lut (.A(\buffer[3] [5]), .B(\buffer[1] [5]), .C(\sendcount[1] ), 
         .Z(n32328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22880_else_3_lut.init = 16'hcaca;
    FD1S3IX select__i7 (.D(n15625), .CK(debug_c_c), .CD(n34073), .Q(\select[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i7.GSR = "ENABLED";
    FD1S3IX select__i5 (.D(n32123), .CK(debug_c_c), .CD(n34073), .Q(\select[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i5.GSR = "ENABLED";
    FD1S3IX select__i4 (.D(n32122), .CK(debug_c_c), .CD(n34073), .Q(\select[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i4.GSR = "ENABLED";
    FD1S3IX select__i3 (.D(n32121), .CK(debug_c_c), .CD(n34073), .Q(\select[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i3.GSR = "ENABLED";
    FD1S3IX select__i2 (.D(n15641), .CK(debug_c_c), .CD(n34073), .Q(\select[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i2.GSR = "ENABLED";
    FD1S3IX select__i1 (.D(n32120), .CK(debug_c_c), .CD(n34073), .Q(\select[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i1.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i31 (.D(\buffer[5] [7]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i31.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i30 (.D(\buffer[5] [6]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i30.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i29 (.D(\buffer[5] [5]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i29.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i28 (.D(\buffer[5] [4]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i28.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i3 (.D(n9241[3]), .SP(n13567), .CD(n16519), .CK(debug_c_c), 
            .Q(esc_data[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i3.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i27 (.D(\buffer[5] [3]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i27.GSR = "ENABLED";
    LUT4 mux_1564_i16_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[15]), 
         .D(n224_adj_56[15]), .Z(n3948[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i16_3_lut_4_lut.init = 16'hf780;
    FD1P3AX databus_out_i0_i26 (.D(\buffer[5] [2]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i26.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i25 (.D(\buffer[5] [1]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i25.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i24 (.D(\buffer[5] [0]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i24.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i23 (.D(\buffer[4] [7]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i23.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i22 (.D(\buffer[4] [6]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i22.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i21 (.D(\buffer[4] [5]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i21.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i20 (.D(\buffer[4] [4]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i20.GSR = "ENABLED";
    LUT4 i4_2_lut_rep_454 (.A(n1432), .B(n1414[15]), .Z(n32275)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_2_lut_rep_454.init = 16'heeee;
    FD1P3IX esc_data_i0_i5 (.D(n9241[5]), .SP(n13567), .CD(n16519), .CK(debug_c_c), 
            .Q(esc_data[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i5.GSR = "ENABLED";
    LUT4 i23334_then_3_lut (.A(\buffer[0] [0]), .B(\buffer[2] [0]), .C(\sendcount[1] ), 
         .Z(n32332)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23334_then_3_lut.init = 16'hcaca;
    LUT4 i23334_else_3_lut (.A(\buffer[3] [0]), .B(\buffer[1] [0]), .C(\sendcount[1] ), 
         .Z(n32331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23334_else_3_lut.init = 16'hcaca;
    FD1P3AX databus_out_i0_i19 (.D(\buffer[4] [3]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i19.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i18 (.D(\buffer[4] [2]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i18.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i17 (.D(\buffer[4] [1]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i17.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i16 (.D(\buffer[4] [0]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i16.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i15 (.D(\buffer[3] [7]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i15.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i6 (.D(n9241[6]), .SP(n13567), .CD(n16519), .CK(debug_c_c), 
            .Q(esc_data[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i6.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i14 (.D(\buffer[3] [6]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i14.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i13 (.D(\buffer[3] [5]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i13.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i12 (.D(\buffer[3] [4]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i12.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i11 (.D(\buffer[3] [3]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i11.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i10 (.D(\buffer[3] [2]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i10.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i7 (.D(n9241[7]), .SP(n13567), .CD(n16519), .CK(debug_c_c), 
            .Q(esc_data[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i7.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i9 (.D(\buffer[3] [1]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i9.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i8 (.D(\buffer[3] [0]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i8.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i7 (.D(\buffer[2] [7]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i7.GSR = "ENABLED";
    LUT4 mux_1564_i15_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[14]), 
         .D(n224_adj_56[14]), .Z(n3948[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i15_3_lut_4_lut.init = 16'hf780;
    FD1P3AX databus_out_i0_i6 (.D(\buffer[2] [6]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i6.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i5 (.D(\buffer[2] [5]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i5.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i4 (.D(\buffer[2] [4]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i4.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i3 (.D(\buffer[2] [3]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i3.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i2 (.D(\buffer[2] [2]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i2.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i1 (.D(\buffer[2] [1]), .SP(n2748), .CK(debug_c_c), 
            .Q(databus_out[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i1.GSR = "ENABLED";
    LUT4 mux_1564_i14_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[13]), 
         .D(n224_adj_56[13]), .Z(n3948[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_408_3_lut (.A(n1432), .B(n1414[15]), .C(n1414[12]), 
         .Z(n32229)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_408_3_lut.init = 16'hfefe;
    FD1P3AX esc_data_i0_i4 (.D(n5765[4]), .SP(n13567), .CK(debug_c_c), 
            .Q(esc_data[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i4.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i2 (.D(n5765[2]), .SP(n13567), .CK(debug_c_c), 
            .Q(esc_data[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i2.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i1 (.D(n5765[1]), .SP(n13567), .CK(debug_c_c), 
            .Q(esc_data[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i1.GSR = "ENABLED";
    LUT4 mux_1564_i13_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[12]), 
         .D(n224_adj_56[12]), .Z(n3948[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i13_3_lut_4_lut.init = 16'hf780;
    FD1S3IX bufcount__i3 (.D(n32321), .CK(debug_c_c), .CD(n34073), .Q(bufcount[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i3.GSR = "ENABLED";
    FD1S3IX bufcount__i2 (.D(n34061), .CK(debug_c_c), .CD(n34073), .Q(bufcount[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i2.GSR = "ENABLED";
    FD1S3IX bufcount__i1 (.D(n15654), .CK(debug_c_c), .CD(n34073), .Q(bufcount[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i1.GSR = "ENABLED";
    LUT4 i22883_then_3_lut (.A(\buffer[0] [4]), .B(\buffer[2] [4]), .C(\sendcount[1] ), 
         .Z(n32335)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22883_then_3_lut.init = 16'hcaca;
    LUT4 i22883_else_3_lut (.A(\buffer[3] [4]), .B(\buffer[1] [4]), .C(\sendcount[1] ), 
         .Z(n32334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22883_else_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_455 (.A(n1414[19]), .B(n1414[3]), .C(n1414[11]), 
         .Z(n32276)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_455.init = 16'hfefe;
    LUT4 i15842_3_lut_rep_356 (.A(n1414[13]), .B(n32213), .C(n1432), .Z(n32177)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i15842_3_lut_rep_356.init = 16'hc8c8;
    LUT4 mux_1564_i12_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[11]), 
         .D(n224_adj_56[11]), .Z(n3948[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i12_3_lut_4_lut.init = 16'hf780;
    FD1P3AX tx_data_i0_i4 (.D(n2156[4]), .SP(n32180), .CK(debug_c_c), 
            .Q(tx_data[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n2156[3]), .SP(n32180), .CK(debug_c_c), 
            .Q(tx_data[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i1 (.D(n2156[1]), .SP(n32180), .CK(debug_c_c), 
            .Q(tx_data[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    LUT4 i22886_then_3_lut (.A(\buffer[0] [3]), .B(\buffer[2] [3]), .C(\sendcount[1] ), 
         .Z(n32338)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22886_then_3_lut.init = 16'hcaca;
    LUT4 i22886_else_3_lut (.A(\buffer[3] [3]), .B(\buffer[1] [3]), .C(\sendcount[1] ), 
         .Z(n32337)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22886_else_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i11_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[10]), 
         .D(n224_adj_56[10]), .Z(n3948[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i22889_then_3_lut (.A(\buffer[0] [2]), .B(\buffer[2] [2]), .C(\sendcount[1] ), 
         .Z(n32341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22889_then_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i10_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[9]), 
         .D(n224_adj_56[9]), .Z(n3948[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 i22889_else_3_lut (.A(\buffer[3] [2]), .B(\buffer[1] [2]), .C(\sendcount[1] ), 
         .Z(n32340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22889_else_3_lut.init = 16'hcaca;
    LUT4 mux_1564_i9_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[8]), 
         .D(n224_adj_56[8]), .Z(n3948[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 i22895_then_3_lut (.A(\buffer[0] [1]), .B(\buffer[2] [1]), .C(\sendcount[1] ), 
         .Z(n32344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22895_then_3_lut.init = 16'hcaca;
    LUT4 i22895_else_3_lut (.A(\buffer[3] [1]), .B(\buffer[1] [1]), .C(\sendcount[1] ), 
         .Z(n32343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22895_else_3_lut.init = 16'hcaca;
    LUT4 i22874_then_3_lut (.A(\buffer[0] [7]), .B(\buffer[2] [7]), .C(\sendcount[1] ), 
         .Z(n32347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22874_then_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_53 (.A(n32172), .B(n32278), .C(n34065), 
         .D(register_addr[0]), .Z(n13545)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_53.init = 16'hf4f0;
    LUT4 i22874_else_3_lut (.A(\buffer[3] [7]), .B(\buffer[1] [7]), .C(\sendcount[1] ), 
         .Z(n32346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22874_else_3_lut.init = 16'hcaca;
    LUT4 i3_2_lut_4_lut (.A(n1414[19]), .B(n1414[3]), .C(n1414[11]), .D(n29532), 
         .Z(n9_adj_38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_2_lut_4_lut.init = 16'hfffe;
    LUT4 n29702_bdd_4_lut (.A(bufcount[1]), .B(n1414[4]), .C(bufcount[0]), 
         .D(bufcount[3]), .Z(n32397)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam n29702_bdd_4_lut.init = 16'h0080;
    LUT4 n29702_bdd_4_lut_23775 (.A(n29702), .B(n32280), .C(n1414[0]), 
         .D(n1414[3]), .Z(n32395)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C)) */ ;
    defparam n29702_bdd_4_lut_23775.init = 16'hdd0f;
    LUT4 mux_1564_i8_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[7]), 
         .D(n224_adj_56[7]), .Z(n3948[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1564_i7_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[6]), 
         .D(n224_adj_56[6]), .Z(n3948[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1564_i6_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[5]), 
         .D(n224_adj_56[5]), .Z(n3948[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1564_i5_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[4]), 
         .D(n224_adj_56[4]), .Z(n3948[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1564_i4_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[3]), 
         .D(n224_adj_56[3]), .Z(n3948[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_457 (.A(\select[2] ), .B(prev_select), .Z(n32278)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_457.init = 16'h2222;
    LUT4 mux_1564_i3_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[2]), 
         .D(n224_adj_56[2]), .Z(n3948[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut (.A(n1414[3]), .B(n29702), .C(n1414[13]), .Z(n14_c)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut.init = 16'hf2f2;
    LUT4 i1_2_lut_2_lut_3_lut (.A(\select[2] ), .B(prev_select), .C(n34065), 
         .Z(n2760)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_2_lut_3_lut.init = 16'h0202;
    LUT4 i1_2_lut_3_lut_adj_54 (.A(n1414[3]), .B(n29702), .C(\buffer[2] [0]), 
         .Z(n29720)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_54.init = 16'h2020;
    LUT4 mux_1564_i2_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[1]), 
         .D(n224_adj_56[1]), .Z(n3948[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_adj_55 (.A(n1414[3]), .B(n29702), .C(\buffer[2] [1]), 
         .Z(n29727)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_55.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_56 (.A(n1414[3]), .B(n29702), .C(\buffer[2] [2]), 
         .Z(n29721)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_56.init = 16'h2020;
    LUT4 i1_2_lut_rep_458 (.A(register_addr[5]), .B(register_addr[4]), .Z(n32279)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_458.init = 16'heeee;
    LUT4 i1_2_lut_4_lut (.A(n29750), .B(rw), .C(n32154), .D(n34065), 
         .Z(n13885)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut.init = 16'hff20;
    LUT4 i1_2_lut_3_lut_adj_57 (.A(n1414[3]), .B(n29702), .C(\buffer[2] [3]), 
         .Z(n29725)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_57.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_58 (.A(n1414[3]), .B(n29702), .C(\buffer[2] [4]), 
         .Z(n29723)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_58.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_59 (.A(n1414[3]), .B(n29702), .C(\buffer[2] [5]), 
         .Z(n29719)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_59.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_60 (.A(n1414[3]), .B(n29702), .C(\buffer[2] [6]), 
         .Z(n29728)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_60.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_61 (.A(n1414[3]), .B(n29702), .C(\buffer[2] [7]), 
         .Z(n29726)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_61.init = 16'h2020;
    LUT4 i23076_2_lut_2_lut_3_lut_4_lut (.A(register_addr[5]), .B(register_addr[4]), 
         .C(n32235), .D(n32315), .Z(n21718)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i23076_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_adj_62 (.A(n1414[3]), .B(n29702), .C(\buffer[3] [0]), 
         .Z(n29724)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_62.init = 16'h2020;
    LUT4 i913_2_lut_rep_459 (.A(escape), .B(debug_c_7), .Z(n32280)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i913_2_lut_rep_459.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_adj_63 (.A(n1414[3]), .B(n29702), .C(\buffer[3] [1]), 
         .Z(n29722)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_63.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_64 (.A(n1414[3]), .B(n29702), .C(\buffer[3] [2]), 
         .Z(n29731)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_64.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_65 (.A(n1414[3]), .B(n29702), .C(\buffer[3] [3]), 
         .Z(n29729)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_65.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_66 (.A(n1414[3]), .B(n29702), .C(\buffer[3] [4]), 
         .Z(n29735)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_66.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_67 (.A(n1414[3]), .B(n29702), .C(\buffer[3] [5]), 
         .Z(n29732)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_67.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_68 (.A(n1414[3]), .B(n29702), .C(\buffer[3] [6]), 
         .Z(n29715)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_68.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_69 (.A(n1414[3]), .B(n29702), .C(\buffer[3] [7]), 
         .Z(n29730)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_69.init = 16'h2020;
    LUT4 i2_3_lut_rep_380_4_lut (.A(escape), .B(debug_c_7), .C(n29702), 
         .D(n1414[4]), .Z(n32201)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i2_3_lut_rep_380_4_lut.init = 16'hffbf;
    LUT4 i1_2_lut_3_lut_adj_70 (.A(n1414[3]), .B(n29702), .C(\buffer[4] [0]), 
         .Z(n29733)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_70.init = 16'h2020;
    LUT4 i1_3_lut_rep_460 (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .Z(n32281)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i1_3_lut_rep_460.init = 16'hecec;
    LUT4 i1_2_lut_3_lut_adj_71 (.A(n1414[3]), .B(n29702), .C(\buffer[4] [1]), 
         .Z(n29716)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_71.init = 16'h2020;
    LUT4 i2_2_lut_rep_409_4_lut (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1414[4]), .Z(n32230)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+!(D))) */ ;
    defparam i2_2_lut_rep_409_4_lut.init = 16'hecff;
    LUT4 i1_2_lut_4_lut_adj_72 (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1414[4]), .Z(n7)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i1_2_lut_4_lut_adj_72.init = 16'hec00;
    LUT4 i1_2_lut_3_lut_adj_73 (.A(n1414[3]), .B(n29702), .C(\buffer[4] [2]), 
         .Z(n29739)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_73.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_74 (.A(n1414[3]), .B(n29702), .C(\buffer[4] [3]), 
         .Z(n29737)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_74.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_75 (.A(n1414[3]), .B(n29702), .C(\buffer[4] [4]), 
         .Z(n29736)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_75.init = 16'h2020;
    LUT4 i132_2_lut_rep_461 (.A(register_addr[2]), .B(register_addr[3]), 
         .Z(n32282)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i132_2_lut_rep_461.init = 16'heeee;
    LUT4 i23103_3_lut_4_lut (.A(n32177), .B(n1432), .C(sendcount[4]), 
         .D(n30294), .Z(n14_adj_39)) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A (C (D)+!C !(D)))) */ ;
    defparam i23103_3_lut_4_lut.init = 16'h0dd0;
    LUT4 i2_2_lut_rep_412_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[4]), .D(register_addr[5]), .Z(n32233)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_2_lut_rep_412_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_76 (.A(n1414[3]), .B(n29702), .C(\buffer[4] [5]), 
         .Z(n29734)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_76.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_77 (.A(n1414[3]), .B(n29702), .C(\buffer[4] [6]), 
         .Z(n29742)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_77.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_78 (.A(n1414[3]), .B(n29702), .C(\buffer[4] [7]), 
         .Z(n29741)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_78.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_79 (.A(n1414[3]), .B(n29702), .C(\buffer[5] [0]), 
         .Z(n29738)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_79.init = 16'h2020;
    LUT4 i15550_2_lut_rep_414_3_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[1]), .Z(n32235)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i15550_2_lut_rep_414_3_lut.init = 16'hfefe;
    LUT4 n32395_bdd_4_lut (.A(n32395), .B(n1414[4]), .C(n32397), .D(bufcount[2]), 
         .Z(n34061)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n32395_bdd_4_lut.init = 16'heef0;
    LUT4 i1_2_lut_3_lut_adj_80 (.A(n1414[3]), .B(n29702), .C(\buffer[5] [1]), 
         .Z(n29745)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_80.init = 16'h2020;
    LUT4 mux_1542_i18_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[17]), 
         .D(n224[17]), .Z(n3862[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_adj_81 (.A(n1414[3]), .B(n29702), .C(\buffer[5] [2]), 
         .Z(n29740)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_81.init = 16'h2020;
    LUT4 i23143_2_lut_rep_381_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[0]), .D(register_addr[1]), .Z(n32202)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i23143_2_lut_rep_381_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_rep_410_3_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[1]), .Z(n32231)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_rep_410_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_adj_82 (.A(n1414[3]), .B(n29702), .C(\buffer[5] [3]), 
         .Z(n29743)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_82.init = 16'h2020;
    LUT4 i2_3_lut_rep_316_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(n29750), .D(n29983), .Z(n32137)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_3_lut_rep_316_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_adj_83 (.A(n1414[3]), .B(n29702), .C(\buffer[5] [4]), 
         .Z(n29744)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_83.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_84 (.A(n1414[3]), .B(n29702), .C(\buffer[5] [5]), 
         .Z(n29717)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_84.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_85 (.A(n1414[3]), .B(n29702), .C(\buffer[5] [6]), 
         .Z(n29746)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_85.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_86 (.A(n1414[3]), .B(n29702), .C(\buffer[5] [7]), 
         .Z(n29718)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_86.init = 16'h2020;
    FD1P3AX send_491 (.D(n12484), .SP(n28225), .CK(debug_c_c), .Q(send));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam send_491.GSR = "ENABLED";
    LUT4 mux_1542_i16_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[15]), 
         .D(n224[15]), .Z(n3862[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_468 (.A(esc_data[5]), .B(esc_data[6]), .Z(n32289)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_468.init = 16'heeee;
    LUT4 n31812_bdd_2_lut_3_lut (.A(esc_data[5]), .B(esc_data[6]), .C(n31812), 
         .Z(n31813)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam n31812_bdd_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_adj_87 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n30052)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_87.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_88 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n30053)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_88.init = 16'hbfbf;
    LUT4 equal_190_i4_2_lut_rep_470 (.A(bufcount[1]), .B(bufcount[2]), .Z(n32291)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam equal_190_i4_2_lut_rep_470.init = 16'heeee;
    PFUMX i8904 (.BLUT(n15624), .ALUT(n28639), .C0(n1867), .Z(n15625));
    LUT4 i2856_2_lut_rep_418_3_lut (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[3]), 
         .Z(n32239)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i2856_2_lut_rep_418_3_lut.init = 16'hfefe;
    LUT4 mux_1542_i1_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[0]), 
         .D(n224[0]), .Z(n3862[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_adj_89 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n30023)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_89.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_90 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n30022)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_90.init = 16'hbfbf;
    LUT4 mux_1542_i15_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[14]), 
         .D(n224[14]), .Z(n3862[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_471 (.A(n1432), .B(sendcount[4]), .Z(n32292)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_471.init = 16'h2222;
    LUT4 n1_bdd_2_lut_23608_3_lut (.A(n1432), .B(sendcount[4]), .C(n31814), 
         .Z(n31815)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam n1_bdd_2_lut_23608_3_lut.init = 16'h2020;
    LUT4 i23105_3_lut_4_lut (.A(\buffer[0] [2]), .B(n29547), .C(\buffer[0] [0]), 
         .D(\buffer[0] [1]), .Z(n28639)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i23105_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_91 (.A(\buffer[0] [2]), .B(n29547), .C(\buffer[0] [1]), 
         .Z(n30012)) /* synthesis lut_function=((B+(C))+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i1_2_lut_3_lut_adj_91.init = 16'hfdfd;
    LUT4 i1_2_lut_3_lut_adj_92 (.A(\buffer[0] [2]), .B(n29547), .C(\buffer[0] [0]), 
         .Z(n30083)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i1_2_lut_3_lut_adj_92.init = 16'hefef;
    LUT4 i23115_3_lut_4_lut (.A(\buffer[0] [2]), .B(n29547), .C(\buffer[0] [1]), 
         .D(\buffer[0] [0]), .Z(n28299)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i23115_3_lut_4_lut.init = 16'h0010;
    LUT4 i23067_4_lut (.A(n32253), .B(n32279), .C(n112), .D(register_addr[2]), 
         .Z(n30075)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;
    defparam i23067_4_lut.init = 16'h0111;
    LUT4 n31121_bdd_3_lut_4_lut (.A(sendcount[2]), .B(n32268), .C(n32333), 
         .D(n31121), .Z(n31122)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam n31121_bdd_3_lut_4_lut.init = 16'hf960;
    LUT4 mux_1542_i14_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[13]), 
         .D(n224[13]), .Z(n3862[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_429_Mux_1_i7_4_lut_4_lut (.A(n32269), .B(n32223), .C(n4_c), 
         .D(n32345), .Z(n9241[1])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_1_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_2_i7_4_lut_4_lut (.A(n32269), .B(n32223), .C(n4_adj_44), 
         .D(n32342), .Z(n9241[2])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_2_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_4_i7_4_lut_4_lut (.A(n32269), .B(n32223), .C(n4_adj_45), 
         .D(n32336), .Z(n9241[4])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_4_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_7_i7_4_lut_4_lut (.A(n32269), .B(n32223), .C(n4_adj_46), 
         .D(n32348), .Z(n9241[7])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_7_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_6_i7_4_lut_4_lut (.A(n32269), .B(n32223), .C(n4_adj_47), 
         .D(n32327), .Z(n9241[6])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_6_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_5_i7_4_lut_4_lut (.A(n32269), .B(n32223), .C(n4_adj_48), 
         .D(n32330), .Z(n9241[5])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_5_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 reduce_or_451_i1_3_lut_4_lut (.A(n32239), .B(n13115), .C(\buffer[0] [7]), 
         .D(n1414[9]), .Z(n1519)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(158[15] 160[18])
    defparam reduce_or_451_i1_3_lut_4_lut.init = 16'hff80;
    LUT4 mux_429_Mux_3_i7_4_lut_4_lut (.A(n32269), .B(n32223), .C(n4_adj_49), 
         .D(n32339), .Z(n9241[3])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_3_i7_4_lut_4_lut.init = 16'hdc10;
    PFUMX i8920 (.BLUT(n15640), .ALUT(n28299), .C0(n1867), .Z(n15641));
    LUT4 i5_3_lut_4_lut (.A(n1414[12]), .B(n32275), .C(n10), .D(n1414[13]), 
         .Z(debug_c_5)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(n1414[4]), .B(n32281), .C(bufcount[0]), 
         .D(n32201), .Z(n28238)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'hd222;
    LUT4 mux_1542_i13_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[12]), 
         .D(n224[12]), .Z(n3862[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1542_i12_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[11]), 
         .D(n224[11]), .Z(n3862[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_93 (.A(n32239), .B(debug_c_7), .C(n13115), .D(n8), 
         .Z(n29368)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_93.init = 16'hdc50;
    LUT4 i1_3_lut (.A(n15), .B(n1414[1]), .C(n1414[0]), .Z(n8)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut.init = 16'hecec;
    LUT4 i4_4_lut (.A(rx_data[2]), .B(n29707), .C(rx_data[5]), .D(n6_adj_52), 
         .Z(n13115)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i4_4_lut.init = 16'h0800;
    LUT4 i2_4_lut_adj_94 (.A(escape), .B(n13_c), .C(debug_c_7), .D(n13034), 
         .Z(n29707)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_4_lut_adj_94.init = 16'h1000;
    LUT4 i1_2_lut_adj_95 (.A(n1414[3]), .B(rx_data[0]), .Z(n6_adj_52)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_95.init = 16'h8888;
    LUT4 i20_2_lut_3_lut_4_lut (.A(n32282), .B(n32279), .C(rw), .D(n32251), 
         .Z(n52)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i20_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_360_3_lut_4_lut (.A(n32282), .B(n32279), .C(prev_select_adj_41), 
         .D(n32251), .Z(n32181)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_360_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_484 (.A(register_addr[4]), .B(register_addr[5]), .Z(n32305)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_484.init = 16'h2222;
    LUT4 i14891_2_lut_rep_361_3_lut_4_lut (.A(register_addr[5]), .B(n32315), 
         .C(\select[3] ), .D(register_addr[4]), .Z(n32182)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i14891_2_lut_rep_361_3_lut_4_lut.init = 16'he0f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_96 (.A(register_addr[4]), .B(register_addr[5]), 
         .C(n32235), .D(n32315), .Z(n29713)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_96.init = 16'h0002;
    LUT4 i15103_2_lut_rep_357_3_lut_4_lut (.A(register_addr[5]), .B(n32315), 
         .C(\select[3] ), .D(register_addr[4]), .Z(n32178)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i15103_2_lut_rep_357_3_lut_4_lut.init = 16'h1000;
    LUT4 i3_4_lut (.A(rx_data[4]), .B(rx_data[3]), .C(rx_data[1]), .D(n29552), 
         .Z(n15)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_97 (.A(n1414[4]), .B(debug_c_7), .C(n1414[2]), .D(n29645), 
         .Z(n29276)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_97.init = 16'heeea;
    LUT4 i1_4_lut_adj_98 (.A(n15), .B(n1414[3]), .C(n1414[0]), .D(n30328), 
         .Z(n29645)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (C+!(D))+!B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_98.init = 16'h50dc;
    LUT4 i15098_2_lut (.A(bufcount[0]), .B(n1414[0]), .Z(n15359)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i15098_2_lut.init = 16'h2222;
    LUT4 i22825_3_lut (.A(n12924), .B(escape), .C(n15), .Z(n30328)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i22825_3_lut.init = 16'hecec;
    LUT4 i24_3_lut_4_lut (.A(bufcount[0]), .B(n32291), .C(rx_data[0]), 
         .D(\buffer[0] [0]), .Z(n11)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_99 (.A(bufcount[0]), .B(n32291), .C(rx_data[1]), 
         .D(\buffer[0] [1]), .Z(n11_adj_54)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_99.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_100 (.A(bufcount[0]), .B(n32291), .C(\buffer[0] [2]), 
         .D(rx_data[2]), .Z(n11_adj_55)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_100.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_101 (.A(bufcount[0]), .B(n32291), .C(\buffer[0] [3]), 
         .D(rx_data[3]), .Z(n11_adj_56)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_101.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_102 (.A(bufcount[0]), .B(n32291), .C(rx_data[4]), 
         .D(\buffer[0] [4]), .Z(n11_adj_57)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_102.init = 16'hfe10;
    LUT4 i5210_3_lut (.A(debug_c_7), .B(n1414[3]), .C(n1414[2]), .Z(n11928)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5210_3_lut.init = 16'h5454;
    LUT4 i23125_3_lut (.A(debug_c_7), .B(n29575), .C(n1414[3]), .Z(n29634)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i23125_3_lut.init = 16'h2020;
    LUT4 i3_4_lut_adj_103 (.A(n30284), .B(n31805), .C(rx_data[0]), .D(escape), 
         .Z(n29575)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_103.init = 16'h0040;
    LUT4 i24_3_lut_4_lut_adj_104 (.A(bufcount[0]), .B(n32291), .C(\buffer[0] [5]), 
         .D(rx_data[5]), .Z(n11_adj_58)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_104.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_105 (.A(bufcount[0]), .B(n32291), .C(\buffer[0] [6]), 
         .D(rx_data[6]), .Z(n11_adj_59)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_105.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_106 (.A(bufcount[0]), .B(n32291), .C(\buffer[0] [7]), 
         .D(rx_data[7]), .Z(n11_adj_60)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_106.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_107 (.A(bufcount[0]), .B(n32291), .C(\buffer[1] [0]), 
         .D(rx_data[0]), .Z(n11_adj_61)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_107.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_108 (.A(bufcount[0]), .B(n32291), .C(\buffer[1] [1]), 
         .D(rx_data[1]), .Z(n11_adj_62)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_108.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_109 (.A(bufcount[0]), .B(n32291), .C(rx_data[2]), 
         .D(\buffer[1] [2]), .Z(n11_adj_63)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_109.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_110 (.A(bufcount[0]), .B(n32291), .C(\buffer[1] [3]), 
         .D(rx_data[3]), .Z(n11_adj_64)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_110.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_111 (.A(bufcount[0]), .B(n32291), .C(\buffer[1] [4]), 
         .D(rx_data[4]), .Z(n11_adj_65)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_111.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_112 (.A(bufcount[0]), .B(n32291), .C(\buffer[1] [5]), 
         .D(rx_data[5]), .Z(n11_adj_66)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_112.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_113 (.A(bufcount[0]), .B(n32291), .C(rx_data[6]), 
         .D(\buffer[1] [6]), .Z(n11_adj_67)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_113.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_114 (.A(bufcount[0]), .B(n32291), .C(rx_data[7]), 
         .D(\buffer[1] [7]), .Z(n11_adj_68)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_114.init = 16'hfd20;
    LUT4 n6_bdd_4_lut (.A(esc_data[3]), .B(esc_data[2]), .C(esc_data[4]), 
         .D(esc_data[1]), .Z(n31812)) /* synthesis lut_function=(A (B+!(C (D)))+!A !(B (C (D))+!B !(C+(D)))) */ ;
    defparam n6_bdd_4_lut.init = 16'h9ffe;
    LUT4 mux_1542_i17_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[16]), 
         .D(n224[16]), .Z(n3862[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1542_i30_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[29]), 
         .D(n224[29]), .Z(n3862[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i30_3_lut_4_lut.init = 16'hf780;
    LUT4 reduce_or_457_i1_3_lut (.A(busy), .B(n1414[13]), .C(n1414[20]), 
         .Z(n1525)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam reduce_or_457_i1_3_lut.init = 16'hdcdc;
    LUT4 i459_2_lut (.A(n5774), .B(n1432), .Z(n1526)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i459_2_lut.init = 16'h4444;
    LUT4 i944_3_lut (.A(n1414[5]), .B(n32213), .C(n1414[10]), .Z(n2746)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i944_3_lut.init = 16'hc8c8;
    LUT4 i1_2_lut_3_lut_adj_115 (.A(rx_data[1]), .B(rx_data[4]), .C(rx_data[3]), 
         .Z(n13034)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i1_2_lut_3_lut_adj_115.init = 16'h0808;
    LUT4 i1_2_lut_rep_493 (.A(register_addr[5]), .B(register_addr[4]), .Z(n32314)) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_493.init = 16'hdddd;
    LUT4 i23131_3_lut_3_lut_4_lut (.A(register_addr[5]), .B(register_addr[4]), 
         .C(n32235), .D(n32315), .Z(n28302)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i23131_3_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i4442_3_lut (.A(n1414[16]), .B(n2687), .C(busy), .Z(n11158)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4442_3_lut.init = 16'hcece;
    LUT4 i5211_3_lut (.A(busy), .B(n1414[17]), .C(n1414[16]), .Z(n11930)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5211_3_lut.init = 16'ha8a8;
    LUT4 i1_2_lut_3_lut_4_lut_adj_116 (.A(n32291), .B(bufcount[3]), .C(\buffer[0] [7]), 
         .D(n13115), .Z(n29924)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_116.init = 16'h0e00;
    LUT4 n12742_bdd_2_lut_23725 (.A(sendcount[0]), .B(sendcount[3]), .Z(n31117)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam n12742_bdd_2_lut_23725.init = 16'hbbbb;
    LUT4 i2_4_lut_adj_117 (.A(n35), .B(busy), .C(n31815), .D(n1414[17]), 
         .Z(n29278)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_117.init = 16'hfbfa;
    LUT4 mux_1542_i11_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[10]), 
         .D(n224[10]), .Z(n3862[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_118 (.A(n1414[15]), .B(esc_data[7]), .C(n31813), 
         .D(esc_data[0]), .Z(n35)) /* synthesis lut_function=(A (B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_118.init = 16'ha8aa;
    LUT4 mux_1542_i10_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[9]), 
         .D(n224[9]), .Z(n3862[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1542_i9_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[8]), 
         .D(n224[8]), .Z(n3862[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 i4435_3_lut (.A(n1414[19]), .B(n1414[18]), .C(busy), .Z(n11151)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4435_3_lut.init = 16'hcece;
    LUT4 i5212_3_lut (.A(busy), .B(n1414[20]), .C(n1414[19]), .Z(n11932)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5212_3_lut.init = 16'ha8a8;
    LUT4 i1_4_lut_adj_119 (.A(n1414[4]), .B(\buffer[0] [1]), .C(n11_adj_54), 
         .D(n14_c), .Z(n29244)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_119.init = 16'heca0;
    LUT4 i1_4_lut_adj_120 (.A(n1414[4]), .B(\buffer[0] [2]), .C(n11_adj_55), 
         .D(n14_c), .Z(n29204)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_120.init = 16'heca0;
    FD1S3AX escape_501 (.D(n10915), .CK(debug_c_c), .Q(escape));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam escape_501.GSR = "ENABLED";
    FD1P3AX rw_498 (.D(n1414[10]), .SP(n2746), .CK(debug_c_c), .Q(rw));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_121 (.A(n1414[4]), .B(\buffer[0] [3]), .C(n11_adj_56), 
         .D(n14_c), .Z(n29202)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_121.init = 16'heca0;
    PFUMX i23737 (.BLUT(n32319), .ALUT(n32320), .C0(n32201), .Z(n32321));
    LUT4 i1_4_lut_adj_122 (.A(n1414[4]), .B(\buffer[0] [4]), .C(n11_adj_57), 
         .D(n14_c), .Z(n29218)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_122.init = 16'heca0;
    LUT4 i1_4_lut_adj_123 (.A(n1414[4]), .B(\buffer[0] [5]), .C(n11_adj_58), 
         .D(n14_c), .Z(n29208)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_123.init = 16'heca0;
    LUT4 i23060_2_lut_rep_335_3_lut (.A(n1414[13]), .B(n32213), .C(n1432), 
         .Z(n32156)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i23060_2_lut_rep_335_3_lut.init = 16'h0808;
    LUT4 i2_4_lut_adj_124 (.A(databus[17]), .B(n5), .C(n1414[13]), .D(n29716), 
         .Z(n28156)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_124.init = 16'hffec;
    LUT4 i1_4_lut_adj_125 (.A(n29903), .B(debug_c_7), .C(n1414[0]), .D(n1414[1]), 
         .Z(n13422)) /* synthesis lut_function=(A+!(B+!(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_125.init = 16'hbbba;
    LUT4 i1_4_lut_adj_126 (.A(n1414[4]), .B(\buffer[0] [6]), .C(n11_adj_59), 
         .D(n14_c), .Z(n29200)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_126.init = 16'heca0;
    LUT4 i3_4_lut_adj_127 (.A(sendcount[3]), .B(n32268), .C(sendcount[2]), 
         .D(n32292), .Z(n29903)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_127.init = 16'h0200;
    LUT4 i1_4_lut_adj_128 (.A(n1414[4]), .B(\buffer[0] [7]), .C(n11_adj_60), 
         .D(n14_c), .Z(n29214)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_128.init = 16'heca0;
    LUT4 i1_4_lut_adj_129 (.A(n1414[4]), .B(\buffer[1] [0]), .C(n11_adj_61), 
         .D(n14_c), .Z(n29210)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_129.init = 16'heca0;
    LUT4 i2_3_lut_rep_495 (.A(register_addr[3]), .B(register_addr[4]), .C(register_addr[2]), 
         .Z(n32316)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_495.init = 16'hfefe;
    LUT4 i1_4_lut_adj_130 (.A(n1414[4]), .B(\buffer[1] [1]), .C(n11_adj_62), 
         .D(n14_c), .Z(n29224)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_130.init = 16'heca0;
    LUT4 i1_2_lut_rep_431_4_lut (.A(register_addr[3]), .B(register_addr[4]), 
         .C(register_addr[2]), .D(register_addr[5]), .Z(n32252)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_431_4_lut.init = 16'h0100;
    LUT4 i1_4_lut_adj_131 (.A(n1414[4]), .B(\buffer[1] [2]), .C(n11_adj_63), 
         .D(n14_c), .Z(n29242)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_131.init = 16'heca0;
    LUT4 i1_4_lut_adj_132 (.A(n1414[4]), .B(\buffer[1] [3]), .C(n11_adj_64), 
         .D(n14_c), .Z(n29216)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_132.init = 16'heca0;
    LUT4 i1_4_lut_adj_133 (.A(n1414[4]), .B(\buffer[1] [4]), .C(n11_adj_65), 
         .D(n14_c), .Z(n29220)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_133.init = 16'heca0;
    LUT4 i1_4_lut_adj_134 (.A(n1414[4]), .B(\buffer[0] [0]), .C(n11), 
         .D(n14_c), .Z(n29226)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_134.init = 16'heca0;
    LUT4 i1_4_lut_adj_135 (.A(n1414[4]), .B(\buffer[1] [5]), .C(n11_adj_66), 
         .D(n14_c), .Z(n29222)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_135.init = 16'heca0;
    LUT4 i1_4_lut_adj_136 (.A(n1414[4]), .B(\buffer[1] [6]), .C(n11_adj_67), 
         .D(n14_c), .Z(n29228)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_136.init = 16'heca0;
    LUT4 i1_4_lut_adj_137 (.A(n1414[4]), .B(\buffer[1] [7]), .C(n11_adj_68), 
         .D(n14_c), .Z(n29230)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_137.init = 16'heca0;
    LUT4 i23040_4_lut (.A(n7), .B(n30316), .C(n32280), .D(n1414[3]), 
         .Z(n9411)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C+!(D))))) */ ;
    defparam i23040_4_lut.init = 16'h0544;
    LUT4 i2_4_lut_adj_138 (.A(databus[0]), .B(n5_adj_73), .C(n1414[13]), 
         .D(n29720), .Z(n28134)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_138.init = 16'hffec;
    LUT4 select_2118_Select_16_i5_4_lut (.A(\buffer[2] [0]), .B(n1414[4]), 
         .C(rx_data[0]), .D(n30023), .Z(n5_adj_73)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_16_i5_4_lut.init = 16'h88c0;
    LUT4 i22813_3_lut (.A(n1414[13]), .B(n1414[0]), .C(n1414[4]), .Z(n30316)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22813_3_lut.init = 16'hfefe;
    LUT4 i2_4_lut_adj_139 (.A(databus[1]), .B(n5_adj_74), .C(n1414[13]), 
         .D(n29727), .Z(n28136)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_139.init = 16'hffec;
    LUT4 select_2118_Select_17_i5_4_lut (.A(\buffer[2] [1]), .B(n1414[4]), 
         .C(rx_data[1]), .D(n30023), .Z(n5_adj_74)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_17_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_140 (.A(databus[2]), .B(n5_adj_75), .C(n1414[13]), 
         .D(n29721), .Z(n28104)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_140.init = 16'hffec;
    LUT4 select_2118_Select_18_i5_4_lut (.A(\buffer[2] [2]), .B(n1414[4]), 
         .C(rx_data[2]), .D(n30023), .Z(n5_adj_75)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_18_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_141 (.A(databus[3]), .B(n5_adj_76), .C(n1414[13]), 
         .D(n29725), .Z(n28106)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_141.init = 16'hffec;
    LUT4 select_2118_Select_19_i5_4_lut (.A(\buffer[2] [3]), .B(n1414[4]), 
         .C(rx_data[3]), .D(n30023), .Z(n5_adj_76)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_19_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_142 (.A(databus[4]), .B(n5_adj_77), .C(n1414[13]), 
         .D(n29723), .Z(n28137)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_142.init = 16'hffec;
    LUT4 select_2118_Select_20_i5_4_lut (.A(\buffer[2] [4]), .B(n1414[4]), 
         .C(rx_data[4]), .D(n30023), .Z(n5_adj_77)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_20_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_143 (.A(databus[5]), .B(n5_adj_78), .C(n1414[13]), 
         .D(n29719), .Z(n28143)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_143.init = 16'hffec;
    LUT4 select_2118_Select_21_i5_4_lut (.A(\buffer[2] [5]), .B(n1414[4]), 
         .C(rx_data[5]), .D(n30023), .Z(n5_adj_78)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_21_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_144 (.A(databus[6]), .B(n5_adj_79), .C(n1414[13]), 
         .D(n29728), .Z(n28147)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_144.init = 16'hffec;
    LUT4 select_2118_Select_22_i5_4_lut (.A(\buffer[2] [6]), .B(n1414[4]), 
         .C(rx_data[6]), .D(n30023), .Z(n5_adj_79)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_22_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_145 (.A(databus[7]), .B(n5_adj_80), .C(n1414[13]), 
         .D(n29726), .Z(n28145)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_145.init = 16'hffec;
    LUT4 select_2118_Select_23_i5_4_lut (.A(\buffer[2] [7]), .B(n1414[4]), 
         .C(rx_data[7]), .D(n30023), .Z(n5_adj_80)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_23_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_146 (.A(databus[8]), .B(n5_adj_81), .C(n1414[13]), 
         .D(n29724), .Z(n28146)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_146.init = 16'hffec;
    LUT4 select_2118_Select_24_i5_4_lut (.A(\buffer[3] [0]), .B(n1414[4]), 
         .C(rx_data[0]), .D(n30022), .Z(n5_adj_81)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_24_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_147 (.A(databus[9]), .B(n5_adj_82), .C(n1414[13]), 
         .D(n29722), .Z(n28142)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_147.init = 16'hffec;
    LUT4 i1_2_lut_adj_148 (.A(n34065), .B(n13576), .Z(n13899)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_148.init = 16'heeee;
    LUT4 select_2118_Select_25_i5_4_lut (.A(\buffer[3] [1]), .B(n1414[4]), 
         .C(rx_data[1]), .D(n30022), .Z(n5_adj_82)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_25_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_149 (.A(databus[10]), .B(n5_adj_83), .C(n1414[13]), 
         .D(n29731), .Z(n28149)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_149.init = 16'hffec;
    LUT4 select_2118_Select_26_i5_4_lut (.A(\buffer[3] [2]), .B(n1414[4]), 
         .C(rx_data[2]), .D(n30022), .Z(n5_adj_83)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_26_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_150 (.A(databus[11]), .B(n5_adj_84), .C(n1414[13]), 
         .D(n29729), .Z(n28153)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_150.init = 16'hffec;
    LUT4 select_2118_Select_27_i5_4_lut (.A(\buffer[3] [3]), .B(n1414[4]), 
         .C(rx_data[3]), .D(n30022), .Z(n5_adj_84)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_27_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_151 (.A(databus[12]), .B(n5_adj_85), .C(n1414[13]), 
         .D(n29735), .Z(n28150)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_151.init = 16'hffec;
    LUT4 select_2118_Select_28_i5_4_lut (.A(\buffer[3] [4]), .B(n1414[4]), 
         .C(rx_data[4]), .D(n30022), .Z(n5_adj_85)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_28_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_152 (.A(databus[13]), .B(n5_adj_86), .C(n1414[13]), 
         .D(n29732), .Z(n28152)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_152.init = 16'hffec;
    LUT4 select_2118_Select_29_i5_4_lut (.A(\buffer[3] [5]), .B(n1414[4]), 
         .C(rx_data[5]), .D(n30022), .Z(n5_adj_86)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_29_i5_4_lut.init = 16'h88c0;
    LUT4 i3341_2_lut_3_lut_4_lut_4_lut (.A(bufcount[1]), .B(n32201), .C(n32230), 
         .D(bufcount[0]), .Z(n1810[1])) /* synthesis lut_function=(A (B (C+!(D)))+!A !((C+!(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i3341_2_lut_3_lut_4_lut_4_lut.init = 16'h8488;
    LUT4 i2_4_lut_adj_153 (.A(databus[14]), .B(n5_adj_87), .C(n1414[13]), 
         .D(n29715), .Z(n28151)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_153.init = 16'hffec;
    LUT4 select_2118_Select_30_i5_4_lut (.A(\buffer[3] [6]), .B(n1414[4]), 
         .C(rx_data[6]), .D(n30022), .Z(n5_adj_87)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_30_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_4_lut_adj_154 (.A(n32252), .B(n32165), .C(n29750), .D(n34065), 
         .Z(n13769)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_4_lut_adj_154.init = 16'hff80;
    LUT4 i2_4_lut_adj_155 (.A(databus[15]), .B(n5_adj_88), .C(n1414[13]), 
         .D(n29730), .Z(n28148)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_155.init = 16'hffec;
    LUT4 i1_2_lut_adj_156 (.A(register_addr[0]), .B(\control_reg[7] ), .Z(n8585)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_156.init = 16'h4444;
    LUT4 i1_2_lut_rep_347_3_lut_4_lut (.A(register_addr[3]), .B(n32315), 
         .C(\select[4] ), .D(register_addr[2]), .Z(n32168)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_347_3_lut_4_lut.init = 16'h0010;
    LUT4 i15399_2_lut_3_lut (.A(n1414[0]), .B(n1414[8]), .C(\select[1] ), 
         .Z(n15661)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i15399_2_lut_3_lut.init = 16'h1010;
    LUT4 i15137_2_lut_3_lut (.A(n1414[0]), .B(n1414[8]), .C(\select[3] ), 
         .Z(n16363)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i15137_2_lut_3_lut.init = 16'h1010;
    LUT4 i15337_2_lut_3_lut (.A(n1414[0]), .B(n1414[8]), .C(\select[7] ), 
         .Z(n15624)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i15337_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_157 (.A(n1414[0]), .B(n1414[8]), .C(\select[4] ), 
         .Z(n16289)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_157.init = 16'h1010;
    LUT4 n29902_bdd_4_lut (.A(sendcount[3]), .B(sendcount[2]), .C(sendcount[0]), 
         .D(\sendcount[1] ), .Z(n31814)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam n29902_bdd_4_lut.init = 16'h4001;
    LUT4 i15336_2_lut_3_lut (.A(n1414[0]), .B(n1414[8]), .C(\select[5] ), 
         .Z(n15626)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i15336_2_lut_3_lut.init = 16'h1010;
    LUT4 rx_data_2__bdd_4_lut (.A(rx_data[2]), .B(rx_data[3]), .C(rx_data[4]), 
         .D(rx_data[1]), .Z(n31805)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D))+!B !(C+(D))))) */ ;
    defparam rx_data_2__bdd_4_lut.init = 16'h6001;
    LUT4 select_2118_Select_31_i5_4_lut (.A(\buffer[3] [7]), .B(n1414[4]), 
         .C(rx_data[7]), .D(n30022), .Z(n5_adj_88)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_31_i5_4_lut.init = 16'h88c0;
    LUT4 i15393_2_lut_3_lut (.A(n1414[0]), .B(n1414[8]), .C(\select[2] ), 
         .Z(n15640)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i15393_2_lut_3_lut.init = 16'h1010;
    LUT4 select_2118_Select_33_i5_4_lut (.A(\buffer[4] [1]), .B(n1414[4]), 
         .C(rx_data[1]), .D(n30052), .Z(n5)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_33_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_158 (.A(databus[16]), .B(n5_adj_89), .C(n1414[13]), 
         .D(n29733), .Z(n28154)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_158.init = 16'hffec;
    LUT4 i2_3_lut_rep_319_4_lut (.A(prev_select_adj_42), .B(n32163), .C(rw), 
         .D(n29750), .Z(n32140)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_319_4_lut.init = 16'h0400;
    LUT4 select_2118_Select_32_i5_4_lut (.A(\buffer[4] [0]), .B(n1414[4]), 
         .C(rx_data[0]), .D(n30052), .Z(n5_adj_89)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_32_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_159 (.A(databus[18]), .B(n5_adj_91), .C(n1414[13]), 
         .D(n29739), .Z(n28157)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_159.init = 16'hffec;
    LUT4 i2_3_lut_4_lut (.A(prev_select_adj_42), .B(n32163), .C(n13118), 
         .D(n29977), .Z(n4034)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut.init = 16'h4000;
    LUT4 select_2118_Select_34_i5_4_lut (.A(\buffer[4] [2]), .B(n1414[4]), 
         .C(rx_data[2]), .D(n30052), .Z(n5_adj_91)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_34_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_160 (.A(databus[19]), .B(n5_adj_92), .C(n1414[13]), 
         .D(n29737), .Z(n28161)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_160.init = 16'hffec;
    LUT4 mux_1542_i29_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[28]), 
         .D(n224[28]), .Z(n3862[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i29_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1542_i28_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[27]), 
         .D(n224[27]), .Z(n3862[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i28_3_lut_4_lut.init = 16'hf780;
    LUT4 select_2118_Select_35_i5_4_lut (.A(\buffer[4] [3]), .B(n1414[4]), 
         .C(rx_data[3]), .D(n30052), .Z(n5_adj_92)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_35_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_161 (.A(databus[20]), .B(n5_adj_93), .C(n1414[13]), 
         .D(n29736), .Z(n28105)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_161.init = 16'hffec;
    LUT4 select_2118_Select_36_i5_4_lut (.A(\buffer[4] [4]), .B(n1414[4]), 
         .C(rx_data[4]), .D(n30052), .Z(n5_adj_93)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_36_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_162 (.A(databus[21]), .B(n5_adj_94), .C(n1414[13]), 
         .D(n29734), .Z(n28172)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_162.init = 16'hffec;
    LUT4 select_2118_Select_37_i5_4_lut (.A(\buffer[4] [5]), .B(n1414[4]), 
         .C(rx_data[5]), .D(n30052), .Z(n5_adj_94)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_37_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_163 (.A(databus[22]), .B(n5_adj_95), .C(n1414[13]), 
         .D(n29742), .Z(n28162)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_163.init = 16'hffec;
    LUT4 select_2118_Select_38_i5_4_lut (.A(\buffer[4] [6]), .B(n1414[4]), 
         .C(rx_data[6]), .D(n30052), .Z(n5_adj_95)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_38_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_164 (.A(databus[23]), .B(n5_adj_96), .C(n1414[13]), 
         .D(n29741), .Z(n28168)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_164.init = 16'hffec;
    LUT4 mux_1884_i3_3_lut (.A(n9241[2]), .B(sendcount[0]), .C(n5774), 
         .Z(n5765[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1884_i3_3_lut.init = 16'hcaca;
    LUT4 select_2118_Select_39_i5_4_lut (.A(\buffer[4] [7]), .B(n1414[4]), 
         .C(rx_data[7]), .D(n30052), .Z(n5_adj_96)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_39_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_165 (.A(databus[24]), .B(n5_adj_97), .C(n1414[13]), 
         .D(n29738), .Z(n28163)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_165.init = 16'hffec;
    LUT4 select_2118_Select_40_i5_4_lut (.A(\buffer[5] [0]), .B(n1414[4]), 
         .C(rx_data[0]), .D(n30053), .Z(n5_adj_97)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_40_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_166 (.A(databus[25]), .B(n5_adj_98), .C(n1414[13]), 
         .D(n29745), .Z(n28169)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_166.init = 16'hffec;
    LUT4 mux_1564_i24_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[23]), 
         .D(n224_adj_56[23]), .Z(n3948[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 select_2118_Select_41_i5_4_lut (.A(\buffer[5] [1]), .B(n1414[4]), 
         .C(rx_data[1]), .D(n30053), .Z(n5_adj_98)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_41_i5_4_lut.init = 16'h88c0;
    LUT4 i15844_3_lut_rep_359 (.A(n2687), .B(n32213), .C(n1414[18]), .Z(n32180)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i15844_3_lut_rep_359.init = 16'hc8c8;
    LUT4 i2_4_lut_adj_167 (.A(databus[26]), .B(n5_adj_100), .C(n1414[13]), 
         .D(n29740), .Z(n28165)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_167.init = 16'hffec;
    LUT4 select_2118_Select_42_i5_4_lut (.A(\buffer[5] [2]), .B(n1414[4]), 
         .C(rx_data[2]), .D(n30053), .Z(n5_adj_100)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_42_i5_4_lut.init = 16'h88c0;
    LUT4 mux_429_Mux_2_i4_3_lut (.A(\buffer[4] [2]), .B(\buffer[5] [2]), 
         .C(sendcount[0]), .Z(n4_adj_44)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_2_i4_3_lut.init = 16'hacac;
    LUT4 i23089_2_lut_3_lut (.A(n2687), .B(n32213), .C(n1414[18]), .Z(n16522)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i23089_2_lut_3_lut.init = 16'h0808;
    LUT4 i2_4_lut_adj_168 (.A(databus[27]), .B(n5_adj_101), .C(n1414[13]), 
         .D(n29743), .Z(n28171)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_168.init = 16'hffec;
    LUT4 i1_2_lut_adj_169 (.A(rw), .B(\select[2] ), .Z(n64)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_169.init = 16'h8888;
    LUT4 select_2118_Select_43_i5_4_lut (.A(\buffer[5] [3]), .B(n1414[4]), 
         .C(rx_data[3]), .D(n30053), .Z(n5_adj_101)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_43_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_adj_170 (.A(n1414[6]), .B(n1414[11]), .Z(n1867)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_170.init = 16'heeee;
    LUT4 i1_2_lut_adj_171 (.A(register_addr[0]), .B(\control_reg[7]_adj_43 ), 
         .Z(n8594)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_171.init = 16'h4444;
    LUT4 i2_4_lut_adj_172 (.A(databus[28]), .B(n5_adj_103), .C(n1414[13]), 
         .D(n29744), .Z(n28166)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_172.init = 16'hffec;
    LUT4 select_2118_Select_44_i5_4_lut (.A(\buffer[5] [4]), .B(n1414[4]), 
         .C(rx_data[4]), .D(n30053), .Z(n5_adj_103)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_44_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_173 (.A(databus[29]), .B(n5_adj_104), .C(n1414[13]), 
         .D(n29717), .Z(n28170)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_173.init = 16'hffec;
    LUT4 select_2118_Select_45_i5_4_lut (.A(\buffer[5] [5]), .B(n1414[4]), 
         .C(rx_data[5]), .D(n30053), .Z(n5_adj_104)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_45_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_174 (.A(databus[30]), .B(n5_adj_105), .C(n1414[13]), 
         .D(n29746), .Z(n28167)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_174.init = 16'hffec;
    LUT4 select_2118_Select_46_i5_4_lut (.A(\buffer[5] [6]), .B(n1414[4]), 
         .C(rx_data[6]), .D(n30053), .Z(n5_adj_105)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_46_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_175 (.A(databus[31]), .B(n5_adj_106), .C(n1414[13]), 
         .D(n29718), .Z(n28160)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_175.init = 16'hffec;
    LUT4 i1_4_lut_adj_176 (.A(n1414[15]), .B(n7_adj_107), .C(n32_c), .D(n32289), 
         .Z(n2687)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_176.init = 16'h0080;
    LUT4 select_2118_Select_47_i5_4_lut (.A(\buffer[5] [7]), .B(n1414[4]), 
         .C(rx_data[7]), .D(n30053), .Z(n5_adj_106)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_2118_Select_47_i5_4_lut.init = 16'h88c0;
    LUT4 mux_1542_i8_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[7]), 
         .D(n224[7]), .Z(n3862[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_2_lut_adj_177 (.A(esc_data[7]), .B(esc_data[0]), .Z(n7_adj_107)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_2_lut_adj_177.init = 16'h4444;
    LUT4 i9648_then_4_lut (.A(bufcount[3]), .B(n1414[0]), .C(n1414[3]), 
         .D(n1414[4]), .Z(n32320)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i9648_then_4_lut.init = 16'haaa2;
    LUT4 i9648_else_4_lut (.A(bufcount[3]), .B(n1414[0]), .C(n1414[3]), 
         .D(n1414[4]), .Z(n32319)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i9648_else_4_lut.init = 16'h0002;
    LUT4 mux_1542_i7_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[6]), 
         .D(n224[6]), .Z(n3862[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1542_i6_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[5]), 
         .D(n224[5]), .Z(n3862[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1564_i23_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[22]), 
         .D(n224_adj_56[22]), .Z(n3948[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 i3_4_lut_adj_178 (.A(\buffer[0] [3]), .B(\buffer[0] [5]), .C(\buffer[0] [4]), 
         .D(\buffer[0] [6]), .Z(n29547)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i3_4_lut_adj_178.init = 16'hfffe;
    LUT4 mux_1884_i2_3_lut (.A(n9241[1]), .B(sendcount[0]), .C(n5774), 
         .Z(n5765[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1884_i2_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_1_i4_3_lut (.A(\buffer[4] [1]), .B(\buffer[5] [1]), 
         .C(sendcount[0]), .Z(n4_c)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_1_i4_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_adj_179 (.A(register_addr[0]), .B(\control_reg[7]_adj_44 ), 
         .Z(n1)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_179.init = 16'h4444;
    LUT4 mux_510_i5_3_lut (.A(n2687), .B(esc_data[4]), .C(n1414[18]), 
         .Z(n2156[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_510_i5_3_lut.init = 16'hcaca;
    LUT4 i23043_2_lut (.A(sendcount[0]), .B(n9), .Z(n22501)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i23043_2_lut.init = 16'h7777;
    LUT4 i1_4_lut_adj_180 (.A(sendcount[4]), .B(n1_adj_113), .C(n6_adj_114), 
         .D(n12746), .Z(n9)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i1_4_lut_adj_180.init = 16'hfeff;
    FD1P3AX reg_addr_i0_i7 (.D(\buffer[1] [7]), .SP(n2746), .CK(debug_c_c), 
            .Q(register_addr[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i7.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i6 (.D(\buffer[1] [6]), .SP(n2746), .CK(debug_c_c), 
            .Q(register_addr[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i6.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i5 (.D(\buffer[1] [5]), .SP(n2746), .CK(debug_c_c), 
            .Q(register_addr[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i5.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i4 (.D(\buffer[1] [4]), .SP(n2746), .CK(debug_c_c), 
            .Q(register_addr[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i4.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i3 (.D(\buffer[1] [3]), .SP(n2746), .CK(debug_c_c), 
            .Q(register_addr[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i3.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i2 (.D(\buffer[1] [2]), .SP(n2746), .CK(debug_c_c), 
            .Q(register_addr[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i2.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i1 (.D(\buffer[1] [1]), .SP(n2746), .CK(debug_c_c), 
            .Q(register_addr[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i1.GSR = "ENABLED";
    LUT4 mux_510_i4_3_lut (.A(n2687), .B(esc_data[3]), .C(n1414[18]), 
         .Z(n2156[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_510_i4_3_lut.init = 16'hcaca;
    LUT4 equal_634_i1_4_lut (.A(sendcount[0]), .B(n13), .C(n18), .D(n14), 
         .Z(n1_adj_113)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam equal_634_i1_4_lut.init = 16'h5556;
    LUT4 i1_2_lut_rep_334_3_lut_4_lut (.A(register_addr[2]), .B(n32253), 
         .C(n32261), .D(\select[4] ), .Z(n32155)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_334_3_lut_4_lut.init = 16'h1000;
    LUT4 mux_510_i2_3_lut (.A(n2687), .B(esc_data[1]), .C(n1414[18]), 
         .Z(n2156[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_510_i2_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut (.A(n1414[19]), .B(n1414[16]), .C(n12484), .Z(n28225)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i2_3_lut.init = 16'hefef;
    LUT4 i23163_3_lut (.A(n32213), .B(n1414[20]), .C(n1414[17]), .Z(n12484)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i23163_3_lut.init = 16'h0202;
    LUT4 i2_4_lut_adj_181 (.A(\reg_size[2] ), .B(sendcount[3]), .C(sendcount[2]), 
         .D(n32284), .Z(n6_adj_114)) /* synthesis lut_function=(A (B (C+!(D))+!B ((D)+!C))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i2_4_lut_adj_181.init = 16'he7de;
    FD1S3IX state_FSM_i2 (.D(n29368), .CK(debug_c_c), .CD(n34073), .Q(n1414[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i2.GSR = "ENABLED";
    FD1S3IX state_FSM_i3 (.D(n29276), .CK(debug_c_c), .CD(n34073), .Q(n1414[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i3.GSR = "ENABLED";
    FD1S3IX state_FSM_i4 (.D(n11928), .CK(debug_c_c), .CD(n34073), .Q(n1414[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i4.GSR = "ENABLED";
    FD1S3IX state_FSM_i5 (.D(n29634), .CK(debug_c_c), .CD(n32169), .Q(n1414[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i5.GSR = "ENABLED";
    FD1S3IX state_FSM_i6 (.D(n29924), .CK(debug_c_c), .CD(n32169), .Q(n1414[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i6.GSR = "ENABLED";
    FD1S3IX state_FSM_i7 (.D(n1414[5]), .CK(debug_c_c), .CD(n32169), .Q(n1414[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i7.GSR = "ENABLED";
    FD1S3IX state_FSM_i8 (.D(n1414[6]), .CK(debug_c_c), .CD(n32169), .Q(n1414[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i8.GSR = "ENABLED";
    FD1S3IX state_FSM_i9 (.D(n1414[7]), .CK(debug_c_c), .CD(n32169), .Q(n1414[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i9.GSR = "ENABLED";
    FD1S3IX state_FSM_i10 (.D(n1414[8]), .CK(debug_c_c), .CD(n32169), 
            .Q(n1414[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i10.GSR = "ENABLED";
    FD1S3IX state_FSM_i11 (.D(n1519), .CK(debug_c_c), .CD(n32169), .Q(n1414[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i11.GSR = "ENABLED";
    FD1S3IX state_FSM_i12 (.D(n1414[10]), .CK(debug_c_c), .CD(n32169), 
            .Q(n1414[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i12.GSR = "ENABLED";
    FD1S3IX state_FSM_i13 (.D(n1414[11]), .CK(debug_c_c), .CD(n32169), 
            .Q(n1414[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i13.GSR = "ENABLED";
    FD1S3IX state_FSM_i14 (.D(n1414[12]), .CK(debug_c_c), .CD(n32169), 
            .Q(n1414[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i14.GSR = "ENABLED";
    FD1S3IX state_FSM_i15 (.D(n1525), .CK(debug_c_c), .CD(n32169), .Q(n1432));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i15.GSR = "ENABLED";
    FD1S3IX state_FSM_i16 (.D(n1526), .CK(debug_c_c), .CD(n32169), .Q(n1414[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i16.GSR = "ENABLED";
    FD1S3IX state_FSM_i17 (.D(n11158), .CK(debug_c_c), .CD(n32169), .Q(n1414[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i17.GSR = "ENABLED";
    FD1S3IX state_FSM_i18 (.D(n11930), .CK(debug_c_c), .CD(n32169), .Q(n1414[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i18.GSR = "ENABLED";
    FD1S3IX state_FSM_i19 (.D(n29278), .CK(debug_c_c), .CD(n32169), .Q(n1414[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i19.GSR = "ENABLED";
    FD1S3IX state_FSM_i20 (.D(n11151), .CK(debug_c_c), .CD(n32169), .Q(n1414[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i20.GSR = "ENABLED";
    FD1S3IX state_FSM_i21 (.D(n11932), .CK(debug_c_c), .CD(n32169), .Q(n1414[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i21.GSR = "ENABLED";
    FD1P3IX buffer_0___i2 (.D(n29244), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[0] [1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i2.GSR = "ENABLED";
    FD1P3IX buffer_0___i3 (.D(n29204), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[0] [2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i3.GSR = "ENABLED";
    FD1P3IX buffer_0___i4 (.D(n29202), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[0] [3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i4.GSR = "ENABLED";
    FD1P3IX buffer_0___i5 (.D(n29218), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[0] [4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i5.GSR = "ENABLED";
    FD1P3IX buffer_0___i6 (.D(n29208), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[0] [5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i6.GSR = "ENABLED";
    FD1P3IX buffer_0___i7 (.D(n29200), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[0] [6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i7.GSR = "ENABLED";
    FD1P3IX buffer_0___i8 (.D(n29214), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[0] [7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i8.GSR = "ENABLED";
    FD1P3IX buffer_0___i9 (.D(n29210), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[1] [0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i9.GSR = "ENABLED";
    FD1P3IX buffer_0___i10 (.D(n29224), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[1] [1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i10.GSR = "ENABLED";
    FD1P3IX buffer_0___i11 (.D(n29242), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[1] [2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i11.GSR = "ENABLED";
    FD1P3IX buffer_0___i12 (.D(n29216), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[1] [3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i12.GSR = "ENABLED";
    FD1P3IX buffer_0___i13 (.D(n29220), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[1] [4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i13.GSR = "ENABLED";
    FD1P3IX buffer_0___i14 (.D(n29222), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[1] [5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i14.GSR = "ENABLED";
    FD1P3IX buffer_0___i15 (.D(n29228), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[1] [6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i15.GSR = "ENABLED";
    FD1P3IX buffer_0___i16 (.D(n29230), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[1] [7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i16.GSR = "ENABLED";
    FD1P3IX buffer_0___i17 (.D(n28134), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[2] [0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i17.GSR = "ENABLED";
    FD1P3IX buffer_0___i18 (.D(n28136), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[2] [1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i18.GSR = "ENABLED";
    FD1P3IX buffer_0___i19 (.D(n28104), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[2] [2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i19.GSR = "ENABLED";
    FD1P3IX buffer_0___i20 (.D(n28106), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[2] [3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i20.GSR = "ENABLED";
    FD1P3IX buffer_0___i21 (.D(n28137), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[2] [4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i21.GSR = "ENABLED";
    FD1P3IX buffer_0___i22 (.D(n28143), .SP(n9411), .CD(n32169), .CK(debug_c_c), 
            .Q(\buffer[2] [5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i22.GSR = "ENABLED";
    FD1P3IX buffer_0___i23 (.D(n28147), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[2] [6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i23.GSR = "ENABLED";
    FD1P3IX buffer_0___i24 (.D(n28145), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[2] [7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i24.GSR = "ENABLED";
    FD1P3IX buffer_0___i25 (.D(n28146), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[3] [0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i25.GSR = "ENABLED";
    FD1P3IX buffer_0___i26 (.D(n28142), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[3] [1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i26.GSR = "ENABLED";
    FD1P3IX buffer_0___i27 (.D(n28149), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[3] [2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i27.GSR = "ENABLED";
    FD1P3IX buffer_0___i28 (.D(n28153), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[3] [3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i28.GSR = "ENABLED";
    FD1P3IX buffer_0___i29 (.D(n28150), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[3] [4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i29.GSR = "ENABLED";
    FD1P3IX buffer_0___i30 (.D(n28152), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[3] [5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i30.GSR = "ENABLED";
    FD1P3IX buffer_0___i31 (.D(n28151), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[3] [6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i31.GSR = "ENABLED";
    FD1P3IX buffer_0___i32 (.D(n28148), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[3] [7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i32.GSR = "ENABLED";
    FD1P3IX buffer_0___i33 (.D(n28154), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[4] [0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i33.GSR = "ENABLED";
    FD1P3IX buffer_0___i34 (.D(n28156), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[4] [1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i34.GSR = "ENABLED";
    FD1P3IX buffer_0___i35 (.D(n28157), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[4] [2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i35.GSR = "ENABLED";
    FD1P3IX buffer_0___i36 (.D(n28161), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[4] [3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i36.GSR = "ENABLED";
    FD1P3IX buffer_0___i37 (.D(n28105), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[4] [4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i37.GSR = "ENABLED";
    FD1P3IX buffer_0___i38 (.D(n28172), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[4] [5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i38.GSR = "ENABLED";
    FD1P3IX buffer_0___i39 (.D(n28162), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[4] [6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i39.GSR = "ENABLED";
    FD1P3IX buffer_0___i40 (.D(n28168), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[4] [7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i40.GSR = "ENABLED";
    FD1P3IX buffer_0___i41 (.D(n28163), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[5] [0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i41.GSR = "ENABLED";
    FD1P3IX buffer_0___i42 (.D(n28169), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[5] [1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i42.GSR = "ENABLED";
    FD1P3IX buffer_0___i43 (.D(n28165), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[5] [2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i43.GSR = "ENABLED";
    FD1P3IX buffer_0___i44 (.D(n28171), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[5] [3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i44.GSR = "ENABLED";
    FD1P3IX buffer_0___i45 (.D(n28166), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[5] [4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i45.GSR = "ENABLED";
    FD1P3IX buffer_0___i46 (.D(n28170), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[5] [5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i46.GSR = "ENABLED";
    FD1P3IX buffer_0___i47 (.D(n28167), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[5] [6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i47.GSR = "ENABLED";
    FD1P3IX buffer_0___i48 (.D(n28160), .SP(n9411), .CD(n34073), .CK(debug_c_c), 
            .Q(\buffer[5] [7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i48.GSR = "ENABLED";
    LUT4 mux_1542_i5_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[4]), 
         .D(n224[4]), .Z(n3862[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1542_i4_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[3]), 
         .D(n224[3]), .Z(n3862[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_342_3_lut_4_lut (.A(register_addr[2]), .B(n32253), 
         .C(n32305), .D(\select[4] ), .Z(n32163)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_342_3_lut_4_lut.init = 16'h1000;
    LUT4 i496_2_lut (.A(n1414[3]), .B(n1414[4]), .Z(n1815)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i496_2_lut.init = 16'heeee;
    LUT4 mux_1542_i3_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[2]), 
         .D(n224[2]), .Z(n3862[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1542_i2_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[1]), 
         .D(n224[1]), .Z(n3862[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1564_i1_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[0]), 
         .D(n224_adj_56[0]), .Z(n3948[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1564_i32_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[31]), 
         .D(n224_adj_56[31]), .Z(n3948[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i32_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1564_i31_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[30]), 
         .D(n224_adj_56[30]), .Z(n3948[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i31_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1564_i30_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[29]), 
         .D(n224_adj_56[29]), .Z(n3948[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i30_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1564_i29_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[28]), 
         .D(n224_adj_56[28]), .Z(n3948[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i29_3_lut_4_lut.init = 16'hf780;
    LUT4 i3_4_lut_adj_182 (.A(n30284), .B(rx_data[2]), .C(rx_data[1]), 
         .D(n29701), .Z(n29702)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i3_4_lut_adj_182.init = 16'h0100;
    LUT4 i2_4_lut_adj_183 (.A(n32156), .B(sendcount[3]), .C(n9), .D(n10136), 
         .Z(n27934)) /* synthesis lut_function=(!(A+(B ((D)+!C)+!B !(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_4_lut_adj_183.init = 16'h1040;
    LUT4 i2_3_lut_adj_184 (.A(n28062), .B(\control_reg[7]_adj_44 ), .C(n32285), 
         .Z(n34)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_adj_184.init = 16'h0808;
    LUT4 i2_4_lut_adj_185 (.A(rx_data[4]), .B(rx_data[3]), .C(rx_data[0]), 
         .D(rx_data[1]), .Z(n29701)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_4_lut_adj_185.init = 16'h0010;
    LUT4 i22781_3_lut (.A(rx_data[6]), .B(rx_data[7]), .C(rx_data[5]), 
         .Z(n30284)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22781_3_lut.init = 16'hfefe;
    LUT4 i15348_2_lut (.A(bufcount[1]), .B(n1414[0]), .Z(n15653)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i15348_2_lut.init = 16'h2222;
    LUT4 i23036_2_lut_2_lut (.A(n32213), .B(n9411), .Z(n21572)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i23036_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_adj_186 (.A(register_addr[0]), .B(register_addr[1]), .Z(n112)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(453[13:26])
    defparam i1_2_lut_adj_186.init = 16'heeee;
    LUT4 i2_3_lut_adj_187 (.A(n28053), .B(\control_reg[7] ), .C(n32285), 
         .Z(n32)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_adj_187.init = 16'h0808;
    FD1P3AX rw_498_rep_498 (.D(n1414[10]), .SP(n2746), .CK(debug_c_c), 
            .Q(n34064));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498_rep_498.GSR = "ENABLED";
    LUT4 i1_4_lut_then_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(\sendcount[1] ), 
         .D(sendcount[2]), .Z(n32323)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0001;
    LUT4 i5_4_lut (.A(n9_adj_38), .B(n1414[15]), .C(n8_adj_125), .D(n1414[1]), 
         .Z(debug_c_2)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i5_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_adj_188 (.A(n1414[9]), .B(n1414[17]), .Z(n8_adj_125)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_2_lut_adj_188.init = 16'heeee;
    LUT4 i2_3_lut_adj_189 (.A(n1414[13]), .B(n1414[7]), .C(n1414[5]), 
         .Z(n29532)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_3_lut_adj_189.init = 16'hfefe;
    LUT4 i1_4_lut_adj_190 (.A(n1414[2]), .B(n32275), .C(n8_adj_126), .D(n1414[18]), 
         .Z(debug_c_3)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_190.init = 16'hfffe;
    LUT4 i3_4_lut_adj_191 (.A(n1414[7]), .B(n1414[6]), .C(n32276), .D(n1414[10]), 
         .Z(n8_adj_126)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_191.init = 16'hfffe;
    LUT4 i4_4_lut_adj_192 (.A(n1414[6]), .B(n32229), .C(n29532), .D(n6_adj_127), 
         .Z(debug_c_4)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i4_4_lut_adj_192.init = 16'hfffe;
    LUT4 i1_2_lut_adj_193 (.A(n1414[4]), .B(n1414[20]), .Z(n6_adj_127)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_193.init = 16'heeee;
    LUT4 i4_4_lut_adj_194 (.A(n1414[11]), .B(n1414[10]), .C(n1414[8]), 
         .D(n1414[9]), .Z(n10)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut_adj_194.init = 16'hfffe;
    LUT4 i1_2_lut_adj_195 (.A(register_addr[1]), .B(\steps_reg[5] ), .Z(n14_adj_45)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_195.init = 16'h8888;
    LUT4 i2_3_lut_adj_196 (.A(n28049), .B(\control_reg[7]_adj_46 ), .C(n32285), 
         .Z(n32_adj_47)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_adj_196.init = 16'h0808;
    LUT4 mux_510_i1_3_lut (.A(n2687), .B(esc_data[0]), .C(n1414[18]), 
         .Z(n2156[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_510_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_197 (.A(register_addr[1]), .B(\steps_reg[6] ), .Z(n13_adj_48)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_197.init = 16'h8888;
    LUT4 i1_2_lut_adj_198 (.A(register_addr[1]), .B(\steps_reg[3] ), .Z(n12)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_198.init = 16'h8888;
    LUT4 i1_2_lut_adj_199 (.A(sendcount[0]), .B(sendcount[3]), .Z(n4)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_199.init = 16'h4444;
    LUT4 i2_3_lut_adj_200 (.A(n28061), .B(\control_reg[7]_adj_43 ), .C(n32285), 
         .Z(n32_adj_49)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_adj_200.init = 16'h0808;
    LUT4 i1_2_lut_adj_201 (.A(register_addr[1]), .B(\steps_reg[5]_adj_50 ), 
         .Z(n14_adj_51)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_201.init = 16'h8888;
    FD1P3IX sendcount__i1 (.D(n9281[1]), .SP(n32177), .CD(n32156), .CK(debug_c_c), 
            .Q(\sendcount[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i1.GSR = "ENABLED";
    FD1P3IX sendcount__i2 (.D(n9281[2]), .SP(n32177), .CD(n32156), .CK(debug_c_c), 
            .Q(sendcount[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i2.GSR = "ENABLED";
    LUT4 mux_1564_i26_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[25]), 
         .D(n224_adj_56[25]), .Z(n3948[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i26_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_202 (.A(register_addr[1]), .B(\steps_reg[6]_adj_52 ), 
         .Z(n13_adj_53)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_202.init = 16'h8888;
    LUT4 i2_3_lut_4_lut_adj_203 (.A(n32234), .B(n32316), .C(register_addr[0]), 
         .D(register_addr[1]), .Z(n13412)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_203.init = 16'hfeff;
    LUT4 i1_2_lut_adj_204 (.A(register_addr[1]), .B(\steps_reg[3]_adj_54 ), 
         .Z(n12_adj_55)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_204.init = 16'h8888;
    FD1P3AX sendcount__i3 (.D(n27934), .SP(n32177), .CK(debug_c_c), .Q(sendcount[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i3.GSR = "ENABLED";
    LUT4 mux_1564_i22_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[21]), 
         .D(n224_adj_56[21]), .Z(n3948[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1564_i21_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[20]), 
         .D(n224_adj_56[20]), .Z(n3948[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1542_i31_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[30]), 
         .D(n224[30]), .Z(n3862[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i31_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_205 (.A(n5774), .B(n9547[0]), .C(n32213), .D(n1432), 
         .Z(n16519)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_205.init = 16'h8000;
    LUT4 mux_1542_i32_3_lut_4_lut (.A(n13118), .B(n29983), .C(databus[31]), 
         .D(n224[31]), .Z(n3862[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1542_i32_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_429_Mux_3_i4_3_lut (.A(\buffer[4] [3]), .B(\buffer[5] [3]), 
         .C(sendcount[0]), .Z(n4_adj_49)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_3_i4_3_lut.init = 16'hacac;
    LUT4 mux_429_Mux_5_i4_3_lut (.A(\buffer[4] [5]), .B(\buffer[5] [5]), 
         .C(sendcount[0]), .Z(n4_adj_48)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_5_i4_3_lut.init = 16'hacac;
    LUT4 mux_1564_i28_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[27]), 
         .D(n224_adj_56[27]), .Z(n3948[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i28_3_lut_4_lut.init = 16'hf780;
    LUT4 i14938_2_lut (.A(sendcount[3]), .B(sendcount[0]), .Z(n9547[0])) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i14938_2_lut.init = 16'hdddd;
    LUT4 mux_1564_i27_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[26]), 
         .D(n224_adj_56[26]), .Z(n3948[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i27_3_lut_4_lut.init = 16'hf780;
    LUT4 i946_2_lut (.A(n1414[5]), .B(n32213), .Z(n2748)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i946_2_lut.init = 16'h8888;
    LUT4 mux_429_Mux_6_i4_3_lut (.A(\buffer[4] [6]), .B(\buffer[5] [6]), 
         .C(sendcount[0]), .Z(n4_adj_47)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_6_i4_3_lut.init = 16'hacac;
    LUT4 mux_1564_i25_3_lut_4_lut (.A(n13118), .B(n32153), .C(databus[24]), 
         .D(n224_adj_56[24]), .Z(n3948[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1564_i25_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_429_Mux_7_i4_3_lut (.A(\buffer[4] [7]), .B(\buffer[5] [7]), 
         .C(sendcount[0]), .Z(n4_adj_46)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_7_i4_3_lut.init = 16'hacac;
    PFUMX i23336 (.BLUT(n31122), .ALUT(n31117), .C0(n5774), .Z(n31123));
    PFUMX i23755 (.BLUT(n32346), .ALUT(n32347), .C0(sendcount[0]), .Z(n32348));
    PFUMX i23753 (.BLUT(n32343), .ALUT(n32344), .C0(sendcount[0]), .Z(n32345));
    PFUMX i23751 (.BLUT(n32340), .ALUT(n32341), .C0(sendcount[0]), .Z(n32342));
    PFUMX i23749 (.BLUT(n32337), .ALUT(n32338), .C0(sendcount[0]), .Z(n32339));
    PFUMX i23747 (.BLUT(n32334), .ALUT(n32335), .C0(sendcount[0]), .Z(n32336));
    LUT4 mux_1884_i5_3_lut (.A(n9241[4]), .B(sendcount[0]), .C(n5774), 
         .Z(n5765[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1884_i5_3_lut.init = 16'hcaca;
    FD1P3AX sendcount__i4 (.D(n14_adj_39), .SP(n32177), .CK(debug_c_c), 
            .Q(sendcount[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=493, LSE_RLINE=503 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i4.GSR = "ENABLED";
    PFUMX i23745 (.BLUT(n32331), .ALUT(n32332), .C0(sendcount[0]), .Z(n32333));
    PFUMX i23743 (.BLUT(n32328), .ALUT(n32329), .C0(sendcount[0]), .Z(n32330));
    LUT4 mux_429_Mux_4_i4_3_lut (.A(\buffer[4] [4]), .B(\buffer[5] [4]), 
         .C(sendcount[0]), .Z(n4_adj_45)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_4_i4_3_lut.init = 16'hacac;
    PFUMX i23741 (.BLUT(n32325), .ALUT(n32326), .C0(sendcount[0]), .Z(n32327));
    LUT4 i1_2_lut_adj_206 (.A(register_addr[0]), .B(\control_reg[7]_adj_46 ), 
         .Z(n8576)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_206.init = 16'h4444;
    PFUMX i23739 (.BLUT(n32322), .ALUT(n32323), .C0(sendcount[3]), .Z(n5774));
    \UARTTransmitter(baud_div=12)  uart_output (.n32169(n32169), .tx_data({tx_data}), 
            .n32213(n32213), .send(send), .busy(busy), .n34073(n34073), 
            .\reset_count[14] (\reset_count[14] ), .\reset_count[13] (\reset_count[13] ), 
            .\reset_count[12] (\reset_count[12] ), .n29954(n29954), .uart_tx_c(uart_tx_c), 
            .debug_c_c(debug_c_c), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(65[30] 70[52])
    \UARTReceiver(baud_div=12)  uart_input (.debug_c_c(debug_c_c), .n32213(n32213), 
            .rx_data({rx_data}), .n32169(n32169), .uart_rx_c(uart_rx_c), 
            .debug_c_7(debug_c_7), .n34073(n34073), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(60[27] 64[39])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=12) 
//

module \UARTTransmitter(baud_div=12)  (n32169, tx_data, n32213, send, 
            busy, n34073, \reset_count[14] , \reset_count[13] , \reset_count[12] , 
            n29954, uart_tx_c, debug_c_c, GND_net) /* synthesis syn_module_defined=1 */ ;
    output n32169;
    input [7:0]tx_data;
    output n32213;
    input send;
    output busy;
    output n34073;
    input \reset_count[14] ;
    input \reset_count[13] ;
    input \reset_count[12] ;
    input n29954;
    output uart_tx_c;
    input debug_c_c;
    input GND_net;
    
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [3:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n31486;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n9391, n2743, n31898, n17, n30610, n31084, n31085, n103, 
        n7, n10, n104, n21890, n29956, n2, n30374, n32176, n29906, 
        n31484, n31485, n29907, n14621, n30372, n30373;
    
    FD1S3IX state__i0 (.D(n31486), .CK(bclk), .CD(n32169), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n9391), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    LUT4 n2742_bdd_4_lut (.A(n32213), .B(state[3]), .C(n2743), .D(state[2]), 
         .Z(n31898)) /* synthesis lut_function=(!((B (D)+!B !(C (D)))+!A)) */ ;
    defparam n2742_bdd_4_lut.init = 16'h2088;
    LUT4 i27_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), .D(state[3]), 
         .Z(n17)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B !(C+(D))))) */ ;
    defparam i27_4_lut_4_lut.init = 16'h15fe;
    LUT4 i23208_4_lut_4_lut (.A(state[3]), .B(state[1]), .C(state[0]), 
         .D(send), .Z(n30610)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+(C+(D))))) */ ;
    defparam i23208_4_lut_4_lut.init = 16'h7ffe;
    LUT4 n31084_bdd_2_lut (.A(n31084), .B(state[2]), .Z(n31085)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n31084_bdd_2_lut.init = 16'h2222;
    FD1P3IX busy_34 (.D(n103), .SP(n31085), .CD(n34073), .CK(bclk), 
            .Q(busy));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam busy_34.GSR = "ENABLED";
    LUT4 i1_4_lut_rep_392 (.A(\reset_count[14] ), .B(\reset_count[13] ), 
         .C(\reset_count[12] ), .D(n29954), .Z(n32213)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i1_4_lut_rep_392.init = 16'heeea;
    LUT4 i58_1_lut_rep_348_4_lut (.A(\reset_count[14] ), .B(\reset_count[13] ), 
         .C(\reset_count[12] ), .D(n29954), .Z(n32169)) /* synthesis lut_function=(!(A+(B (C+(D))))) */ ;
    defparam i58_1_lut_rep_348_4_lut.init = 16'h1115;
    LUT4 state_2__bdd_4_lut_23893 (.A(state[0]), .B(state[3]), .C(state[1]), 
         .D(send), .Z(n31084)) /* synthesis lut_function=(A (B (C))+!A !(B+(C+!(D)))) */ ;
    defparam state_2__bdd_4_lut_23893.init = 16'h8180;
    LUT4 i58_1_lut_rep_507 (.A(\reset_count[14] ), .B(\reset_count[13] ), 
         .C(\reset_count[12] ), .D(n29954), .Z(n34073)) /* synthesis lut_function=(!(A+(B (C+(D))))) */ ;
    defparam i58_1_lut_rep_507.init = 16'h1115;
    PFUMX Mux_22_i15 (.BLUT(n7), .ALUT(n10), .C0(state[3]), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;
    LUT4 i15204_2_lut (.A(state[1]), .B(state[0]), .Z(n21890)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15204_2_lut.init = 16'heeee;
    LUT4 i1_2_lut (.A(state[1]), .B(state[0]), .Z(n2743)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_50 (.A(send), .B(state[3]), .Z(n29956)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_50.init = 16'h2222;
    LUT4 Mux_22_i7_4_lut (.A(n2), .B(n30374), .C(state[2]), .D(state[1]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    LUT4 i1_3_lut_rep_355 (.A(n32213), .B(state[2]), .C(state[3]), .Z(n32176)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i1_3_lut_rep_355.init = 16'h2a2a;
    LUT4 i1_3_lut_4_lut (.A(n32213), .B(state[2]), .C(state[3]), .D(n2743), 
         .Z(n29906)) /* synthesis lut_function=(!((B (C+(D))+!B !(D))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h2208;
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i15577_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i15577_4_lut.init = 16'hfcee;
    LUT4 state_1__bdd_2_lut (.A(state[3]), .B(state[0]), .Z(n31484)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_1__bdd_2_lut.init = 16'h1111;
    LUT4 state_1__bdd_4_lut (.A(state[1]), .B(state[3]), .C(state[0]), 
         .D(send), .Z(n31485)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(B (C)+!B (C+!(D)))) */ ;
    defparam state_1__bdd_4_lut.init = 16'h8f0e;
    LUT4 i8998_1_lut (.A(state[3]), .Z(n103)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i8998_1_lut.init = 16'h5555;
    LUT4 i1_3_lut (.A(state[1]), .B(n32176), .C(state[0]), .Z(n29907)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4848;
    PFUMX i23409 (.BLUT(n31485), .ALUT(n31484), .C0(state[2]), .Z(n31486));
    FD1P3AX state__i3 (.D(n31898), .SP(n14621), .CK(bclk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n9391), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n9391), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n9391), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n9391), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n9391), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n9391), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n9391), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    FD1P3AX state__i2 (.D(n29906), .SP(n14621), .CK(bclk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    FD1P3AX state__i1 (.D(n29907), .SP(n14621), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    PFUMX i22871 (.BLUT(n30372), .ALUT(n30373), .C0(state[1]), .Z(n30374));
    LUT4 i22869_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n30372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22869_3_lut.init = 16'hcaca;
    LUT4 i22870_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n30373)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22870_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(n32213), .B(state[2]), .C(n29956), .D(n21890), 
         .Z(n9391)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0020;
    LUT4 i23210_2_lut_3_lut (.A(n32213), .B(state[2]), .C(n30610), .Z(n14621)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i23210_2_lut_3_lut.init = 16'hfdfd;
    FD1P3JX tx_35 (.D(n104), .SP(n17), .PD(n32169), .CK(bclk), .Q(uart_tx_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    \ClockDividerP(factor=12)  baud_gen (.bclk(bclk), .debug_c_c(debug_c_c), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12) 
//

module \ClockDividerP(factor=12)  (bclk, debug_c_c, GND_net) /* synthesis syn_module_defined=1 */ ;
    output bclk;
    input debug_c_c;
    input GND_net;
    
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n8412, n27358, n27357;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n27356, n27355, n27354, n27353, n27352, n27351, n27350, 
        n27349, n27348, n27347, n27346, n27345, n27344, n27343, 
        n16570;
    wire [31:0]n102;
    
    wire n27678, n27677, n27676, n27675, n27674, n27673, n27672, 
        n27671, n27670, n55, n56, n4, n52, n44, n35, n54, 
        n48, n36, n27669, n27668, n46, n32, n27667, n50, n40, 
        n27666, n27665, n27664, n27663;
    
    FD1S3AX clk_o_14 (.D(n8412), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D sub_2074_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27358), .S0(n8412));
    defparam sub_2074_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2074_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2074_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2074_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27357), .COUT(n27358));
    defparam sub_2074_add_2_32.INIT0 = 16'h5555;
    defparam sub_2074_add_2_32.INIT1 = 16'h5555;
    defparam sub_2074_add_2_32.INJECT1_0 = "NO";
    defparam sub_2074_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27356), .COUT(n27357));
    defparam sub_2074_add_2_30.INIT0 = 16'h5555;
    defparam sub_2074_add_2_30.INIT1 = 16'h5555;
    defparam sub_2074_add_2_30.INJECT1_0 = "NO";
    defparam sub_2074_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27355), .COUT(n27356));
    defparam sub_2074_add_2_28.INIT0 = 16'h5555;
    defparam sub_2074_add_2_28.INIT1 = 16'h5555;
    defparam sub_2074_add_2_28.INJECT1_0 = "NO";
    defparam sub_2074_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27354), .COUT(n27355));
    defparam sub_2074_add_2_26.INIT0 = 16'h5555;
    defparam sub_2074_add_2_26.INIT1 = 16'h5555;
    defparam sub_2074_add_2_26.INJECT1_0 = "NO";
    defparam sub_2074_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27353), .COUT(n27354));
    defparam sub_2074_add_2_24.INIT0 = 16'h5555;
    defparam sub_2074_add_2_24.INIT1 = 16'h5555;
    defparam sub_2074_add_2_24.INJECT1_0 = "NO";
    defparam sub_2074_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27352), .COUT(n27353));
    defparam sub_2074_add_2_22.INIT0 = 16'h5555;
    defparam sub_2074_add_2_22.INIT1 = 16'h5555;
    defparam sub_2074_add_2_22.INJECT1_0 = "NO";
    defparam sub_2074_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27351), .COUT(n27352));
    defparam sub_2074_add_2_20.INIT0 = 16'h5555;
    defparam sub_2074_add_2_20.INIT1 = 16'h5555;
    defparam sub_2074_add_2_20.INJECT1_0 = "NO";
    defparam sub_2074_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27350), .COUT(n27351));
    defparam sub_2074_add_2_18.INIT0 = 16'h5555;
    defparam sub_2074_add_2_18.INIT1 = 16'h5555;
    defparam sub_2074_add_2_18.INJECT1_0 = "NO";
    defparam sub_2074_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27349), .COUT(n27350));
    defparam sub_2074_add_2_16.INIT0 = 16'h5555;
    defparam sub_2074_add_2_16.INIT1 = 16'h5555;
    defparam sub_2074_add_2_16.INJECT1_0 = "NO";
    defparam sub_2074_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27348), .COUT(n27349));
    defparam sub_2074_add_2_14.INIT0 = 16'h5555;
    defparam sub_2074_add_2_14.INIT1 = 16'h5555;
    defparam sub_2074_add_2_14.INJECT1_0 = "NO";
    defparam sub_2074_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27347), .COUT(n27348));
    defparam sub_2074_add_2_12.INIT0 = 16'h5555;
    defparam sub_2074_add_2_12.INIT1 = 16'h5555;
    defparam sub_2074_add_2_12.INJECT1_0 = "NO";
    defparam sub_2074_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27346), .COUT(n27347));
    defparam sub_2074_add_2_10.INIT0 = 16'h5555;
    defparam sub_2074_add_2_10.INIT1 = 16'h5555;
    defparam sub_2074_add_2_10.INJECT1_0 = "NO";
    defparam sub_2074_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27345), .COUT(n27346));
    defparam sub_2074_add_2_8.INIT0 = 16'h5555;
    defparam sub_2074_add_2_8.INIT1 = 16'h5555;
    defparam sub_2074_add_2_8.INJECT1_0 = "NO";
    defparam sub_2074_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27344), .COUT(n27345));
    defparam sub_2074_add_2_6.INIT0 = 16'h5555;
    defparam sub_2074_add_2_6.INIT1 = 16'h5555;
    defparam sub_2074_add_2_6.INJECT1_0 = "NO";
    defparam sub_2074_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27343), .COUT(n27344));
    defparam sub_2074_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2074_add_2_4.INIT1 = 16'h5555;
    defparam sub_2074_add_2_4.INJECT1_0 = "NO";
    defparam sub_2074_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_2074_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27343));
    defparam sub_2074_add_2_2.INIT0 = 16'h0000;
    defparam sub_2074_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2074_add_2_2.INJECT1_0 = "NO";
    defparam sub_2074_add_2_2.INJECT1_1 = "NO";
    FD1S3IX count_2667__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i0.GSR = "ENABLED";
    FD1S3IX count_2667__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i1.GSR = "ENABLED";
    FD1S3IX count_2667__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i2.GSR = "ENABLED";
    FD1S3IX count_2667__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i3.GSR = "ENABLED";
    FD1S3IX count_2667__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i4.GSR = "ENABLED";
    FD1S3IX count_2667__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i5.GSR = "ENABLED";
    FD1S3IX count_2667__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i6.GSR = "ENABLED";
    FD1S3IX count_2667__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i7.GSR = "ENABLED";
    FD1S3IX count_2667__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i8.GSR = "ENABLED";
    FD1S3IX count_2667__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i9.GSR = "ENABLED";
    FD1S3IX count_2667__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i10.GSR = "ENABLED";
    FD1S3IX count_2667__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i11.GSR = "ENABLED";
    FD1S3IX count_2667__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i12.GSR = "ENABLED";
    FD1S3IX count_2667__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i13.GSR = "ENABLED";
    FD1S3IX count_2667__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i14.GSR = "ENABLED";
    FD1S3IX count_2667__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i15.GSR = "ENABLED";
    FD1S3IX count_2667__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i16.GSR = "ENABLED";
    FD1S3IX count_2667__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i17.GSR = "ENABLED";
    FD1S3IX count_2667__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i18.GSR = "ENABLED";
    FD1S3IX count_2667__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i19.GSR = "ENABLED";
    FD1S3IX count_2667__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i20.GSR = "ENABLED";
    FD1S3IX count_2667__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i21.GSR = "ENABLED";
    FD1S3IX count_2667__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i22.GSR = "ENABLED";
    FD1S3IX count_2667__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i23.GSR = "ENABLED";
    FD1S3IX count_2667__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i24.GSR = "ENABLED";
    FD1S3IX count_2667__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i25.GSR = "ENABLED";
    FD1S3IX count_2667__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i26.GSR = "ENABLED";
    FD1S3IX count_2667__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i27.GSR = "ENABLED";
    FD1S3IX count_2667__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i28.GSR = "ENABLED";
    FD1S3IX count_2667__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i29.GSR = "ENABLED";
    FD1S3IX count_2667__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i30.GSR = "ENABLED";
    FD1S3IX count_2667__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n16570), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667__i31.GSR = "ENABLED";
    CCU2D count_2667_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27678), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_33.INIT1 = 16'h0000;
    defparam count_2667_add_4_33.INJECT1_0 = "NO";
    defparam count_2667_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2667_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27677), .COUT(n27678), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2667_add_4_31.INJECT1_0 = "NO";
    defparam count_2667_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2667_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27676), .COUT(n27677), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2667_add_4_29.INJECT1_0 = "NO";
    defparam count_2667_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2667_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27675), .COUT(n27676), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2667_add_4_27.INJECT1_0 = "NO";
    defparam count_2667_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2667_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27674), .COUT(n27675), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2667_add_4_25.INJECT1_0 = "NO";
    defparam count_2667_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2667_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27673), .COUT(n27674), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2667_add_4_23.INJECT1_0 = "NO";
    defparam count_2667_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2667_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27672), .COUT(n27673), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2667_add_4_21.INJECT1_0 = "NO";
    defparam count_2667_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2667_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27671), .COUT(n27672), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2667_add_4_19.INJECT1_0 = "NO";
    defparam count_2667_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2667_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27670), .COUT(n27671), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2667_add_4_17.INJECT1_0 = "NO";
    defparam count_2667_add_4_17.INJECT1_1 = "NO";
    LUT4 i23123_4_lut (.A(n55), .B(count[1]), .C(n56), .D(n4), .Z(n16570)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23123_4_lut.init = 16'h0400;
    LUT4 i26_4_lut (.A(count[14]), .B(n52), .C(n44), .D(count[6]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i27_4_lut (.A(n35), .B(n54), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(count[3]), .B(count[0]), .Z(n4)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    CCU2D count_2667_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27669), .COUT(n27670), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2667_add_4_15.INJECT1_0 = "NO";
    defparam count_2667_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2667_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27668), .COUT(n27669), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2667_add_4_13.INJECT1_0 = "NO";
    defparam count_2667_add_4_13.INJECT1_1 = "NO";
    LUT4 i23_4_lut (.A(count[24]), .B(n46), .C(n32), .D(count[16]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i15_3_lut (.A(count[15]), .B(count[31]), .C(count[5]), .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i17_4_lut (.A(count[26]), .B(count[12]), .C(count[28]), .D(count[18]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[13]), .B(count[22]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(count[20]), .B(count[4]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i6_2_lut.init = 16'heeee;
    CCU2D count_2667_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27667), .COUT(n27668), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2667_add_4_11.INJECT1_0 = "NO";
    defparam count_2667_add_4_11.INJECT1_1 = "NO";
    LUT4 i25_4_lut (.A(count[25]), .B(n50), .C(n40), .D(count[9]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(count[7]), .B(count[19]), .C(count[11]), .D(count[21]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[8]), .B(count[29]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i21_4_lut (.A(count[2]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i11_2_lut (.A(count[10]), .B(count[17]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i11_2_lut.init = 16'heeee;
    CCU2D count_2667_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27666), .COUT(n27667), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2667_add_4_9.INJECT1_0 = "NO";
    defparam count_2667_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2667_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27665), .COUT(n27666), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2667_add_4_7.INJECT1_0 = "NO";
    defparam count_2667_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2667_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27664), .COUT(n27665), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2667_add_4_5.INJECT1_0 = "NO";
    defparam count_2667_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2667_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27663), .COUT(n27664), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2667_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2667_add_4_3.INJECT1_0 = "NO";
    defparam count_2667_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2667_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27663), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2667_add_4_1.INIT0 = 16'hF000;
    defparam count_2667_add_4_1.INIT1 = 16'h0555;
    defparam count_2667_add_4_1.INJECT1_0 = "NO";
    defparam count_2667_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \UARTReceiver(baud_div=12) 
//

module \UARTReceiver(baud_div=12)  (debug_c_c, n32213, rx_data, n32169, 
            uart_rx_c, debug_c_7, n34073, GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n32213;
    output [7:0]rx_data;
    input n32169;
    input uart_rx_c;
    output debug_c_7;
    input n34073;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [7:0]rdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(22[12:17])
    
    wire n9339, n9341;
    wire [5:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    
    wire n29114, baud_reset, n19, n32241, bclk, n32224, n31437, 
        n32270;
    wire [7:0]n78;
    
    wire n13158, n13, n9355, n32304, n32310, n9357, n32303, n30045, 
        n9359, n9361, n30059, n29, n16389, n16390, n9363, n22480, 
        n25, n27, n29028, n32815, n32814, n34060, n9365, n9367, 
        n21, n23, n28712, n19_adj_31, n13131, n19_adj_32, n9369, 
        n9371, n9373, n9375, n9377, n9379, n9381, n32298, n32300, 
        n30077, n32, n21_adj_33, n30130, n25_adj_34, n4, n31436, 
        n32242, n33, n31438;
    wire [5:0]n6;
    
    wire n4_adj_35;
    
    FD1P3AX rdata_i0_i0 (.D(n9339), .SP(n32213), .CK(debug_c_c), .Q(rdata[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i0.GSR = "ENABLED";
    FD1P3AX data_i0_i0 (.D(n9341), .SP(n32213), .CK(debug_c_c), .Q(rx_data[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i0.GSR = "ENABLED";
    FD1S3IX state__i0 (.D(n29114), .CK(debug_c_c), .CD(n32169), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i0.GSR = "ENABLED";
    FD1S3JX baud_reset_52 (.D(n19), .CK(debug_c_c), .PD(n32169), .Q(baud_reset)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam baud_reset_52.GSR = "ENABLED";
    LUT4 n29783_bdd_4_lut (.A(n32241), .B(state[4]), .C(bclk), .D(n32224), 
         .Z(n31437)) /* synthesis lut_function=(!((B (C (D))+!B !(C (D)))+!A)) */ ;
    defparam n29783_bdd_4_lut.init = 16'h2888;
    LUT4 i3480_3_lut_rep_449 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n32270)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i3480_3_lut_rep_449.init = 16'h8080;
    LUT4 i3487_2_lut_rep_403_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(state[3]), .Z(n32224)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3487_2_lut_rep_403_4_lut.init = 16'h8000;
    LUT4 i1_4_lut (.A(n78[1]), .B(rdata[1]), .C(n13158), .D(n13), .Z(n9355)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i4408_4_lut (.A(uart_rx_c), .B(rdata[1]), .C(n32304), .D(n32310), 
         .Z(n78[1])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4408_4_lut.init = 16'hcacc;
    LUT4 i1_4_lut_adj_27 (.A(n78[2]), .B(rdata[2]), .C(n13158), .D(n13), 
         .Z(n9357)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_27.init = 16'heca0;
    LUT4 i4406_4_lut (.A(uart_rx_c), .B(rdata[2]), .C(n32303), .D(n30045), 
         .Z(n78[2])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4406_4_lut.init = 16'hccca;
    LUT4 i1_2_lut (.A(state[3]), .B(state[2]), .Z(n30045)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_28 (.A(n78[3]), .B(rdata[3]), .C(n13158), .D(n13), 
         .Z(n9359)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_28.init = 16'heca0;
    LUT4 i4404_4_lut (.A(uart_rx_c), .B(rdata[3]), .C(n32310), .D(n30045), 
         .Z(n78[3])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4404_4_lut.init = 16'hccac;
    LUT4 i1_4_lut_adj_29 (.A(n78[4]), .B(rdata[4]), .C(n13158), .D(n13), 
         .Z(n9361)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_29.init = 16'heca0;
    LUT4 i4402_4_lut (.A(uart_rx_c), .B(rdata[4]), .C(state[2]), .D(n30059), 
         .Z(n78[4])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4402_4_lut.init = 16'hccca;
    PFUMX i9669 (.BLUT(n29), .ALUT(n16389), .C0(state[0]), .Z(n16390));
    LUT4 i1_4_lut_adj_30 (.A(n78[5]), .B(rdata[5]), .C(n13158), .D(n13), 
         .Z(n9363)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_30.init = 16'heca0;
    LUT4 i4400_4_lut (.A(uart_rx_c), .B(rdata[5]), .C(state[2]), .D(n22480), 
         .Z(n78[5])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4400_4_lut.init = 16'hcacc;
    PFUMX i40 (.BLUT(n25), .ALUT(n27), .C0(state[0]), .Z(n29028));
    LUT4 n32815_bdd_4_lut (.A(n32815), .B(state[5]), .C(n32814), .D(state[0]), 
         .Z(n34060)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C (D))) */ ;
    defparam n32815_bdd_4_lut.init = 16'hf022;
    LUT4 i1_4_lut_adj_31 (.A(n78[6]), .B(rdata[6]), .C(n13158), .D(n13), 
         .Z(n9365)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_31.init = 16'heca0;
    LUT4 i4398_4_lut (.A(uart_rx_c), .B(rdata[6]), .C(state[2]), .D(n30059), 
         .Z(n78[6])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4398_4_lut.init = 16'hccac;
    LUT4 i1_4_lut_adj_32 (.A(n78[7]), .B(rdata[7]), .C(n13158), .D(n13), 
         .Z(n9367)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_32.init = 16'heca0;
    PFUMX i36 (.BLUT(n21), .ALUT(n23), .C0(state[5]), .Z(n28712));
    LUT4 i4396_4_lut (.A(rdata[7]), .B(uart_rx_c), .C(state[2]), .D(n22480), 
         .Z(n78[7])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4396_4_lut.init = 16'hcaaa;
    FD1S3IX drdy_51 (.D(n19_adj_31), .CK(debug_c_c), .CD(n34073), .Q(debug_c_7));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam drdy_51.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_33 (.A(rdata[1]), .B(rx_data[1]), .C(n13131), .D(n19_adj_32), 
         .Z(n9369)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_33.init = 16'heca0;
    LUT4 i1_4_lut_adj_34 (.A(rdata[2]), .B(rx_data[2]), .C(n13131), .D(n19_adj_32), 
         .Z(n9371)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_34.init = 16'heca0;
    LUT4 i1_4_lut_adj_35 (.A(rdata[3]), .B(rx_data[3]), .C(n13131), .D(n19_adj_32), 
         .Z(n9373)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_35.init = 16'heca0;
    LUT4 i1_4_lut_adj_36 (.A(rdata[4]), .B(rx_data[4]), .C(n13131), .D(n19_adj_32), 
         .Z(n9375)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_36.init = 16'heca0;
    LUT4 i1_4_lut_adj_37 (.A(rdata[5]), .B(rx_data[5]), .C(n13131), .D(n19_adj_32), 
         .Z(n9377)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_37.init = 16'heca0;
    LUT4 i1_4_lut_adj_38 (.A(rdata[6]), .B(rx_data[6]), .C(n13131), .D(n19_adj_32), 
         .Z(n9379)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_38.init = 16'heca0;
    LUT4 i1_4_lut_adj_39 (.A(rdata[7]), .B(rx_data[7]), .C(n13131), .D(n19_adj_32), 
         .Z(n9381)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_39.init = 16'heca0;
    LUT4 i1_4_lut_adj_40 (.A(n78[0]), .B(rdata[0]), .C(n13158), .D(n13), 
         .Z(n9339)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_40.init = 16'heca0;
    LUT4 i4448_4_lut (.A(uart_rx_c), .B(rdata[0]), .C(n32304), .D(n32303), 
         .Z(n78[0])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i4448_4_lut.init = 16'hccca;
    LUT4 i2_3_lut (.A(state[0]), .B(state[5]), .C(state[4]), .Z(n13)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_477 (.A(state[1]), .B(state[4]), .Z(n32298)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_477.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[4]), .C(n32300), 
         .D(n32304), .Z(n30077)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_41 (.A(state[1]), .B(state[4]), .C(n32), 
         .D(n32304), .Z(n21_adj_33)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_3_lut_4_lut_adj_41.init = 16'hf0f1;
    LUT4 i22634_2_lut_3_lut_4_lut (.A(state[1]), .B(state[4]), .C(uart_rx_c), 
         .D(n32304), .Z(n30130)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i22634_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_42 (.A(state[1]), .B(state[4]), .C(n32304), 
         .D(state[0]), .Z(n25_adj_34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_3_lut_4_lut_adj_42.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut (.A(state[3]), .B(n32270), .C(state[4]), .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 n29783_bdd_3_lut_4_lut (.A(state[3]), .B(n32270), .C(bclk), .D(state[4]), 
         .Z(n31436)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;
    defparam n29783_bdd_3_lut_4_lut.init = 16'hf708;
    LUT4 state_1__bdd_4_lut (.A(state[1]), .B(n32242), .C(n32), .D(uart_rx_c), 
         .Z(n32815)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+(D))) */ ;
    defparam state_1__bdd_4_lut.init = 16'ha2b3;
    LUT4 i1_4_lut_4_lut (.A(state[3]), .B(n32270), .C(bclk), .D(n32), 
         .Z(n33)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut.init = 16'h6a00;
    LUT4 i9668_3_lut_3_lut (.A(state[3]), .B(n32270), .C(bclk), .Z(n16389)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;
    defparam i9668_3_lut_3_lut.init = 16'ha6a6;
    LUT4 state_1__bdd_2_lut (.A(state[1]), .B(bclk), .Z(n32814)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam state_1__bdd_2_lut.init = 16'h9999;
    LUT4 i14912_2_lut_rep_479 (.A(state[0]), .B(state[5]), .Z(n32300)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14912_2_lut_rep_479.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_43 (.A(state[0]), .B(state[5]), .C(state[4]), 
         .Z(n13158)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_43.init = 16'h1010;
    LUT4 i1_4_lut_adj_44 (.A(rdata[0]), .B(rx_data[0]), .C(n13131), .D(n19_adj_32), 
         .Z(n9341)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_44.init = 16'heca0;
    LUT4 i1_2_lut_rep_482 (.A(state[1]), .B(bclk), .Z(n32303)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i1_2_lut_rep_482.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_adj_45 (.A(state[1]), .B(bclk), .C(state[3]), 
         .Z(n30059)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i1_2_lut_3_lut_adj_45.init = 16'hbfbf;
    LUT4 i2_2_lut_rep_483 (.A(state[3]), .B(state[2]), .Z(n32304)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_2_lut_rep_483.init = 16'heeee;
    LUT4 i1_4_lut_adj_46 (.A(state[4]), .B(state[3]), .C(state[2]), .D(state[1]), 
         .Z(n32)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_46.init = 16'heaaa;
    LUT4 i1_2_lut_rep_421_3_lut_4_lut (.A(state[3]), .B(state[2]), .C(state[4]), 
         .D(state[1]), .Z(n32242)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_421_3_lut_4_lut.init = 16'hfffe;
    LUT4 i15185_2_lut_rep_489 (.A(bclk), .B(state[1]), .Z(n32310)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15185_2_lut_rep_489.init = 16'h8888;
    LUT4 i15794_2_lut_3_lut (.A(bclk), .B(state[1]), .C(state[3]), .Z(n22480)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15794_2_lut_3_lut.init = 16'h8080;
    LUT4 i23083_4_lut (.A(baud_reset), .B(n30077), .C(uart_rx_c), .D(n25_adj_34), 
         .Z(n19)) /* synthesis lut_function=(A (B+(C))+!A !((D)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i23083_4_lut.init = 16'ha8ec;
    LUT4 i1_2_lut_rep_420 (.A(n32), .B(state[5]), .Z(n32241)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_420.init = 16'h2222;
    LUT4 i1_3_lut_4_lut (.A(n32), .B(state[5]), .C(state[0]), .D(bclk), 
         .Z(n29114)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_3_lut_4_lut.init = 16'hf200;
    LUT4 i2_3_lut_4_lut (.A(n32304), .B(n32298), .C(state[0]), .D(state[5]), 
         .Z(n13131)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i2_3_lut_4_lut.init = 16'h0100;
    LUT4 i2_3_lut_4_lut_adj_47 (.A(state[0]), .B(n32298), .C(state[5]), 
         .D(n32304), .Z(n19_adj_32)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_3_lut_4_lut_adj_47.init = 16'hffef;
    LUT4 i23085_4_lut (.A(debug_c_7), .B(n30077), .C(uart_rx_c), .D(n25_adj_34), 
         .Z(n19_adj_31)) /* synthesis lut_function=(A (B+(C))+!A !((D)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i23085_4_lut.init = 16'ha8ec;
    PFUMX i23403 (.BLUT(n31437), .ALUT(n31436), .C0(state[0]), .Z(n31438));
    FD1P3AX rdata_i0_i1 (.D(n9355), .SP(n32213), .CK(debug_c_c), .Q(rdata[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i1.GSR = "ENABLED";
    FD1P3AX rdata_i0_i2 (.D(n9357), .SP(n32213), .CK(debug_c_c), .Q(rdata[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i2.GSR = "ENABLED";
    FD1P3AX rdata_i0_i3 (.D(n9359), .SP(n32213), .CK(debug_c_c), .Q(rdata[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i3.GSR = "ENABLED";
    FD1P3AX rdata_i0_i4 (.D(n9361), .SP(n32213), .CK(debug_c_c), .Q(rdata[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i4.GSR = "ENABLED";
    FD1P3AX rdata_i0_i5 (.D(n9363), .SP(n32213), .CK(debug_c_c), .Q(rdata[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i5.GSR = "ENABLED";
    FD1P3AX rdata_i0_i6 (.D(n9365), .SP(n32213), .CK(debug_c_c), .Q(rdata[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i6.GSR = "ENABLED";
    FD1P3AX rdata_i0_i7 (.D(n9367), .SP(n32213), .CK(debug_c_c), .Q(rdata[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i7.GSR = "ENABLED";
    FD1P3AX data_i0_i1 (.D(n9369), .SP(n32213), .CK(debug_c_c), .Q(rx_data[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i1.GSR = "ENABLED";
    FD1P3AX data_i0_i2 (.D(n9371), .SP(n32213), .CK(debug_c_c), .Q(rx_data[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i2.GSR = "ENABLED";
    FD1P3AX data_i0_i3 (.D(n9373), .SP(n32213), .CK(debug_c_c), .Q(rx_data[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i3.GSR = "ENABLED";
    FD1P3AX data_i0_i4 (.D(n9375), .SP(n32213), .CK(debug_c_c), .Q(rx_data[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i4.GSR = "ENABLED";
    FD1P3AX data_i0_i5 (.D(n9377), .SP(n32213), .CK(debug_c_c), .Q(rx_data[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i5.GSR = "ENABLED";
    FD1P3AX data_i0_i6 (.D(n9379), .SP(n32213), .CK(debug_c_c), .Q(rx_data[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i6.GSR = "ENABLED";
    FD1P3AX data_i0_i7 (.D(n9381), .SP(n32213), .CK(debug_c_c), .Q(rx_data[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i7.GSR = "ENABLED";
    FD1S3IX state__i1 (.D(n34060), .CK(debug_c_c), .CD(n34073), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i1.GSR = "ENABLED";
    FD1S3IX state__i2 (.D(n29028), .CK(debug_c_c), .CD(n34073), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i2.GSR = "ENABLED";
    FD1S3IX state__i3 (.D(n16390), .CK(debug_c_c), .CD(n34073), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i3.GSR = "ENABLED";
    FD1S3IX state__i4 (.D(n31438), .CK(debug_c_c), .CD(n34073), .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i4.GSR = "ENABLED";
    FD1S3IX state__i5 (.D(n28712), .CK(debug_c_c), .CD(n34073), .Q(state[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i5.GSR = "ENABLED";
    LUT4 i22645_4_lut (.A(n6[3]), .B(state[5]), .C(n33), .D(n32242), 
         .Z(n29)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i22645_4_lut.init = 16'h3032;
    LUT4 i14950_2_lut (.A(state[3]), .B(uart_rx_c), .Z(n6[3])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(42[8] 47[12])
    defparam i14950_2_lut.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_48 (.A(state[5]), .B(n30130), .C(state[2]), .D(n21_adj_33), 
         .Z(n25)) /* synthesis lut_function=(!(A+!((C (D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_48.init = 16'h5111;
    LUT4 i41_3_lut (.A(state[1]), .B(state[2]), .C(bclk), .Z(n27)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i41_3_lut.init = 16'hc6c6;
    LUT4 i2_4_lut (.A(bclk), .B(n4), .C(state[0]), .D(n32), .Z(n21)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i2_4_lut.init = 16'h4840;
    LUT4 i38_4_lut (.A(n30130), .B(n32224), .C(state[0]), .D(n4_adj_35), 
         .Z(n23)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i38_4_lut.init = 16'hf535;
    LUT4 i1_2_lut_adj_49 (.A(state[4]), .B(bclk), .Z(n4_adj_35)) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_49.init = 16'hdddd;
    \ClockDividerP(factor=12)_U0  baud_gen (.GND_net(GND_net), .bclk(bclk), 
            .debug_c_c(debug_c_c), .baud_reset(baud_reset)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(25[28] 27[56])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12)_U0 
//

module \ClockDividerP(factor=12)_U0  (GND_net, bclk, debug_c_c, baud_reset) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output bclk;
    input debug_c_c;
    input baud_reset;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27646;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n134;
    
    wire n27645, n27644, n27643, n27642, n27641, n27640, n27639, 
        n27638, n27637, n27636, n27635, n27634, n27633, n27632, 
        n27631, n8377, n2903, n27374, n27373, n27372, n55, n28027, 
        n56, n52, n44, n35, n54, n48, n36, n46, n32, n27371, 
        n50, n40, n27370, n27369, n27368, n27367, n27366, n27365, 
        n27364, n27363, n27362, n27361, n27360, n27359;
    
    CCU2D count_2666_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27646), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_33.INIT1 = 16'h0000;
    defparam count_2666_add_4_33.INJECT1_0 = "NO";
    defparam count_2666_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27645), .COUT(n27646), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2666_add_4_31.INJECT1_0 = "NO";
    defparam count_2666_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27644), .COUT(n27645), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2666_add_4_29.INJECT1_0 = "NO";
    defparam count_2666_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27643), .COUT(n27644), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2666_add_4_27.INJECT1_0 = "NO";
    defparam count_2666_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27642), .COUT(n27643), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2666_add_4_25.INJECT1_0 = "NO";
    defparam count_2666_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27641), .COUT(n27642), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2666_add_4_23.INJECT1_0 = "NO";
    defparam count_2666_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27640), .COUT(n27641), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2666_add_4_21.INJECT1_0 = "NO";
    defparam count_2666_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27639), .COUT(n27640), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2666_add_4_19.INJECT1_0 = "NO";
    defparam count_2666_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27638), .COUT(n27639), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2666_add_4_17.INJECT1_0 = "NO";
    defparam count_2666_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27637), .COUT(n27638), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2666_add_4_15.INJECT1_0 = "NO";
    defparam count_2666_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27636), .COUT(n27637), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2666_add_4_13.INJECT1_0 = "NO";
    defparam count_2666_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27635), .COUT(n27636), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2666_add_4_11.INJECT1_0 = "NO";
    defparam count_2666_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27634), .COUT(n27635), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2666_add_4_9.INJECT1_0 = "NO";
    defparam count_2666_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27633), .COUT(n27634), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2666_add_4_7.INJECT1_0 = "NO";
    defparam count_2666_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27632), .COUT(n27633), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2666_add_4_5.INJECT1_0 = "NO";
    defparam count_2666_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27631), .COUT(n27632), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2666_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2666_add_4_3.INJECT1_0 = "NO";
    defparam count_2666_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2666_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27631), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666_add_4_1.INIT0 = 16'hF000;
    defparam count_2666_add_4_1.INIT1 = 16'h0555;
    defparam count_2666_add_4_1.INJECT1_0 = "NO";
    defparam count_2666_add_4_1.INJECT1_1 = "NO";
    FD1S3IX clk_o_14 (.D(n8377), .CK(debug_c_c), .CD(baud_reset), .Q(bclk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2666__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2903), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i0.GSR = "ENABLED";
    CCU2D sub_2072_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27374), .S0(n8377));
    defparam sub_2072_add_2_cout.INIT0 = 16'h0000;
    defparam sub_2072_add_2_cout.INIT1 = 16'h0000;
    defparam sub_2072_add_2_cout.INJECT1_0 = "NO";
    defparam sub_2072_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27373), .COUT(n27374));
    defparam sub_2072_add_2_32.INIT0 = 16'h5555;
    defparam sub_2072_add_2_32.INIT1 = 16'h5555;
    defparam sub_2072_add_2_32.INJECT1_0 = "NO";
    defparam sub_2072_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27372), .COUT(n27373));
    defparam sub_2072_add_2_30.INIT0 = 16'h5555;
    defparam sub_2072_add_2_30.INIT1 = 16'h5555;
    defparam sub_2072_add_2_30.INJECT1_0 = "NO";
    defparam sub_2072_add_2_30.INJECT1_1 = "NO";
    LUT4 i1101_4_lut (.A(n55), .B(baud_reset), .C(n28027), .D(n56), 
         .Z(n2903)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(23[5] 33[8])
    defparam i1101_4_lut.init = 16'hccdc;
    LUT4 i26_4_lut (.A(count[14]), .B(n52), .C(n44), .D(count[6]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut (.A(count[1]), .B(count[3]), .C(count[0]), .Z(n28027)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i27_4_lut (.A(n35), .B(n54), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i23_4_lut (.A(count[24]), .B(n46), .C(n32), .D(count[16]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i23_4_lut.init = 16'hfffe;
    CCU2D sub_2072_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27371), .COUT(n27372));
    defparam sub_2072_add_2_28.INIT0 = 16'h5555;
    defparam sub_2072_add_2_28.INIT1 = 16'h5555;
    defparam sub_2072_add_2_28.INJECT1_0 = "NO";
    defparam sub_2072_add_2_28.INJECT1_1 = "NO";
    LUT4 i15_3_lut (.A(count[15]), .B(count[31]), .C(count[5]), .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i17_4_lut (.A(count[26]), .B(count[12]), .C(count[28]), .D(count[18]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[13]), .B(count[22]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(count[20]), .B(count[4]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i25_4_lut (.A(count[25]), .B(n50), .C(n40), .D(count[9]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i25_4_lut.init = 16'hfffe;
    CCU2D sub_2072_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27370), .COUT(n27371));
    defparam sub_2072_add_2_26.INIT0 = 16'h5555;
    defparam sub_2072_add_2_26.INIT1 = 16'h5555;
    defparam sub_2072_add_2_26.INJECT1_0 = "NO";
    defparam sub_2072_add_2_26.INJECT1_1 = "NO";
    LUT4 i19_4_lut (.A(count[7]), .B(count[19]), .C(count[11]), .D(count[21]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[8]), .B(count[29]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i21_4_lut (.A(count[2]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i11_2_lut (.A(count[10]), .B(count[17]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_2_lut.init = 16'heeee;
    CCU2D sub_2072_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27369), .COUT(n27370));
    defparam sub_2072_add_2_24.INIT0 = 16'h5555;
    defparam sub_2072_add_2_24.INIT1 = 16'h5555;
    defparam sub_2072_add_2_24.INJECT1_0 = "NO";
    defparam sub_2072_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27368), .COUT(n27369));
    defparam sub_2072_add_2_22.INIT0 = 16'h5555;
    defparam sub_2072_add_2_22.INIT1 = 16'h5555;
    defparam sub_2072_add_2_22.INJECT1_0 = "NO";
    defparam sub_2072_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27367), .COUT(n27368));
    defparam sub_2072_add_2_20.INIT0 = 16'h5555;
    defparam sub_2072_add_2_20.INIT1 = 16'h5555;
    defparam sub_2072_add_2_20.INJECT1_0 = "NO";
    defparam sub_2072_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27366), .COUT(n27367));
    defparam sub_2072_add_2_18.INIT0 = 16'h5555;
    defparam sub_2072_add_2_18.INIT1 = 16'h5555;
    defparam sub_2072_add_2_18.INJECT1_0 = "NO";
    defparam sub_2072_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27365), .COUT(n27366));
    defparam sub_2072_add_2_16.INIT0 = 16'h5555;
    defparam sub_2072_add_2_16.INIT1 = 16'h5555;
    defparam sub_2072_add_2_16.INJECT1_0 = "NO";
    defparam sub_2072_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27364), .COUT(n27365));
    defparam sub_2072_add_2_14.INIT0 = 16'h5555;
    defparam sub_2072_add_2_14.INIT1 = 16'h5555;
    defparam sub_2072_add_2_14.INJECT1_0 = "NO";
    defparam sub_2072_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27363), .COUT(n27364));
    defparam sub_2072_add_2_12.INIT0 = 16'h5555;
    defparam sub_2072_add_2_12.INIT1 = 16'h5555;
    defparam sub_2072_add_2_12.INJECT1_0 = "NO";
    defparam sub_2072_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27362), .COUT(n27363));
    defparam sub_2072_add_2_10.INIT0 = 16'h5555;
    defparam sub_2072_add_2_10.INIT1 = 16'h5555;
    defparam sub_2072_add_2_10.INJECT1_0 = "NO";
    defparam sub_2072_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27361), .COUT(n27362));
    defparam sub_2072_add_2_8.INIT0 = 16'h5555;
    defparam sub_2072_add_2_8.INIT1 = 16'h5555;
    defparam sub_2072_add_2_8.INJECT1_0 = "NO";
    defparam sub_2072_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27360), .COUT(n27361));
    defparam sub_2072_add_2_6.INIT0 = 16'h5555;
    defparam sub_2072_add_2_6.INIT1 = 16'h5555;
    defparam sub_2072_add_2_6.INJECT1_0 = "NO";
    defparam sub_2072_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27359), .COUT(n27360));
    defparam sub_2072_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_2072_add_2_4.INIT1 = 16'h5555;
    defparam sub_2072_add_2_4.INJECT1_0 = "NO";
    defparam sub_2072_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_2072_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27359));
    defparam sub_2072_add_2_2.INIT0 = 16'h0000;
    defparam sub_2072_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_2072_add_2_2.INJECT1_0 = "NO";
    defparam sub_2072_add_2_2.INJECT1_1 = "NO";
    FD1S3IX count_2666__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2903), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i1.GSR = "ENABLED";
    FD1S3IX count_2666__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2903), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i2.GSR = "ENABLED";
    FD1S3IX count_2666__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2903), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i3.GSR = "ENABLED";
    FD1S3IX count_2666__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2903), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i4.GSR = "ENABLED";
    FD1S3IX count_2666__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2903), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i5.GSR = "ENABLED";
    FD1S3IX count_2666__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2903), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i6.GSR = "ENABLED";
    FD1S3IX count_2666__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2903), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i7.GSR = "ENABLED";
    FD1S3IX count_2666__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2903), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i8.GSR = "ENABLED";
    FD1S3IX count_2666__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2903), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i9.GSR = "ENABLED";
    FD1S3IX count_2666__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i10.GSR = "ENABLED";
    FD1S3IX count_2666__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i11.GSR = "ENABLED";
    FD1S3IX count_2666__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i12.GSR = "ENABLED";
    FD1S3IX count_2666__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i13.GSR = "ENABLED";
    FD1S3IX count_2666__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i14.GSR = "ENABLED";
    FD1S3IX count_2666__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i15.GSR = "ENABLED";
    FD1S3IX count_2666__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i16.GSR = "ENABLED";
    FD1S3IX count_2666__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i17.GSR = "ENABLED";
    FD1S3IX count_2666__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i18.GSR = "ENABLED";
    FD1S3IX count_2666__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i19.GSR = "ENABLED";
    FD1S3IX count_2666__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i20.GSR = "ENABLED";
    FD1S3IX count_2666__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i21.GSR = "ENABLED";
    FD1S3IX count_2666__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i22.GSR = "ENABLED";
    FD1S3IX count_2666__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i23.GSR = "ENABLED";
    FD1S3IX count_2666__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i24.GSR = "ENABLED";
    FD1S3IX count_2666__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i25.GSR = "ENABLED";
    FD1S3IX count_2666__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i26.GSR = "ENABLED";
    FD1S3IX count_2666__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i27.GSR = "ENABLED";
    FD1S3IX count_2666__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i28.GSR = "ENABLED";
    FD1S3IX count_2666__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i29.GSR = "ENABLED";
    FD1S3IX count_2666__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i30.GSR = "ENABLED";
    FD1S3IX count_2666__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2903), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2666__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0) 
//

module \ArmPeripheral(axis_haddr=8'b0)  (databus, debug_c_c, n34069, n608, 
            n610, \control_reg[7] , n32149, Stepper_X_En_c, Stepper_X_Dir_c, 
            n13511, Stepper_X_M2_c_2, Stepper_X_M1_c_1, \read_size[2] , 
            n2769, n21617, n34067, n34068, n34071, \read_size[0] , 
            n21718, n34066, Stepper_X_M0_c_0, n579, prev_step_clk, 
            step_clk, prev_select, n32203, read_value, n9485, Stepper_X_Step_c, 
            \register_addr[1] , \register_addr[0] , rw, n32181, n32233, 
            n29750, n32279, n13118, n32231, n32235, n32232, n22529, 
            n14812, n32282, n32314, n32315, n30020, n32305, n28426, 
            n32261, n30019, n32187, limit_c_0, n32159, n34065, n14419, 
            n9478, n1, n34, n28062, VCC_net, GND_net, Stepper_X_nFault_c, 
            n24, n32142) /* synthesis syn_module_defined=1 */ ;
    input [31:0]databus;
    input debug_c_c;
    input n34069;
    input n608;
    input n610;
    output \control_reg[7] ;
    input n32149;
    output Stepper_X_En_c;
    output Stepper_X_Dir_c;
    input n13511;
    output Stepper_X_M2_c_2;
    output Stepper_X_M1_c_1;
    output \read_size[2] ;
    input n2769;
    input n21617;
    input n34067;
    input n34068;
    input n34071;
    output \read_size[0] ;
    input n21718;
    input n34066;
    output Stepper_X_M0_c_0;
    input n579;
    output prev_step_clk;
    output step_clk;
    output prev_select;
    input n32203;
    output [31:0]read_value;
    input n9485;
    output Stepper_X_Step_c;
    input \register_addr[1] ;
    input \register_addr[0] ;
    input rw;
    input n32181;
    input n32233;
    input n29750;
    input n32279;
    input n13118;
    input n32231;
    input n32235;
    input n32232;
    output n22529;
    output n14812;
    input n32282;
    input n32314;
    input n32315;
    output n30020;
    input n32305;
    output n28426;
    input n32261;
    output n30019;
    output n32187;
    input limit_c_0;
    input n32159;
    input n34065;
    input n14419;
    output n9478;
    input n1;
    input n34;
    output n28062;
    input VCC_net;
    input GND_net;
    input Stepper_X_nFault_c;
    input n24;
    input n32142;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]n224;
    
    wire n4121;
    wire [31:0]n4122;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n32150, n13444, n11127;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire limit_latched, n182, prev_limit_latched, n30371, int_step, 
        n30393, n30394, n30395;
    wire [31:0]n100;
    
    wire n1_c, n2, n1_adj_12, n2_adj_13, n1_adj_14, n2_adj_15, n1_adj_16, 
        n2_adj_17, n2_adj_18, n30369, n30370;
    wire [31:0]n6439;
    
    wire fault_latched, n30399, n30400, n30401, n49, n62_adj_21, 
        n58_adj_22, n50_adj_23, n41, n60_adj_24, n54_adj_25, n42_adj_26, 
        n52_adj_27, n38_adj_28, n56_adj_29, n46_adj_30, n27430, n27429, 
        n27428, n27427, n27426, n27425, n27424, n27423, n27422, 
        n27421, n27420, n27419, n27418, n27417, n27416, n27415;
    
    LUT4 mux_1610_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n4121), .Z(n4122[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n4121), 
         .Z(n4122[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i26_3_lut.init = 16'hcaca;
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n32150), .PD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n32150), .PD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n32150), .PD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n32150), .PD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n32150), .PD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n32150), .PD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n32150), .PD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n13444), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n13444), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n32149), .CD(n11127), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n32149), .PD(n34069), 
            .CK(debug_c_c), .Q(Stepper_X_En_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n32149), .PD(n34069), 
            .CK(debug_c_c), .Q(Stepper_X_Dir_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n13511), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n32149), .PD(n34069), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n13511), .CK(debug_c_c), .Q(Stepper_X_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n32149), .PD(n34069), 
            .CK(debug_c_c), .Q(Stepper_X_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    LUT4 mux_1610_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n4121), 
         .Z(n4122[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n4121), 
         .Z(n4122[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i12_3_lut.init = 16'hcaca;
    FD1P3AX read_size__i2 (.D(n21617), .SP(n2769), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n4122[31]), .CK(debug_c_c), .CD(n34067), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n4122[30]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n4122[29]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n4122[28]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n4122[27]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n4122[26]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n4122[0]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n4122[25]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n4122[24]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n4122[23]), .CK(debug_c_c), .CD(n34071), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n4122[22]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n4122[21]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n4122[20]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n4122[19]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n21718), .SP(n2769), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n4122[18]), .CK(debug_c_c), .CD(n34069), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n4122[17]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n4122[16]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n13511), .CK(debug_c_c), .Q(Stepper_X_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n13444), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n32203), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n4122[15]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n4122[14]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n4122[13]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n4122[12]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n4122[11]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n4122[10]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n4122[9]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n4122[8]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n4122[7]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n4122[6]), .CK(debug_c_c), .CD(n34069), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n30371), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n4122[5]), .CK(debug_c_c), .CD(n34069), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n4122[4]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    LUT4 mux_1610_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n4121), 
         .Z(n4122[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n4121), .Z(n4122[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i10_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i3 (.D(n4122[3]), .CK(debug_c_c), .CD(n34067), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n4122[2]), .CK(debug_c_c), .CD(n34067), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n4122[1]), .CK(debug_c_c), .CD(n34067), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 mux_1610_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n4121), .Z(n4122[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n4121), .Z(n4122[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i8_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_X_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    PFUMX i22892 (.BLUT(n30393), .ALUT(n30394), .C0(\register_addr[1] ), 
          .Z(n30395));
    LUT4 i15776_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15776_4_lut.init = 16'hc088;
    LUT4 i15775_4_lut (.A(div_factor_reg[9]), .B(\register_addr[1] ), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15775_4_lut.init = 16'hc088;
    LUT4 i15774_4_lut (.A(div_factor_reg[10]), .B(\register_addr[1] ), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15774_4_lut.init = 16'hc088;
    LUT4 i15773_4_lut (.A(div_factor_reg[11]), .B(\register_addr[1] ), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15773_4_lut.init = 16'hc088;
    LUT4 i15772_4_lut (.A(div_factor_reg[12]), .B(\register_addr[1] ), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15772_4_lut.init = 16'hc088;
    LUT4 i15771_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15771_4_lut.init = 16'hc088;
    LUT4 i15770_4_lut (.A(div_factor_reg[14]), .B(\register_addr[1] ), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15770_4_lut.init = 16'hc088;
    LUT4 i15769_4_lut (.A(div_factor_reg[15]), .B(\register_addr[1] ), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15769_4_lut.init = 16'hc088;
    LUT4 i15768_4_lut (.A(div_factor_reg[16]), .B(\register_addr[1] ), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n100[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15768_4_lut.init = 16'hc088;
    LUT4 i15767_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15767_4_lut.init = 16'hc088;
    LUT4 i15766_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15766_4_lut.init = 16'hc088;
    LUT4 i15765_4_lut (.A(div_factor_reg[19]), .B(\register_addr[1] ), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15765_4_lut.init = 16'hc088;
    LUT4 i15764_4_lut (.A(div_factor_reg[20]), .B(\register_addr[1] ), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n100[20])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15764_4_lut.init = 16'hc088;
    LUT4 i15763_4_lut (.A(div_factor_reg[21]), .B(\register_addr[1] ), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15763_4_lut.init = 16'hc088;
    LUT4 i15762_4_lut (.A(div_factor_reg[22]), .B(\register_addr[1] ), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15762_4_lut.init = 16'hc088;
    LUT4 i15761_4_lut (.A(div_factor_reg[23]), .B(\register_addr[1] ), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n100[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15761_4_lut.init = 16'hc088;
    LUT4 i15760_4_lut (.A(div_factor_reg[24]), .B(\register_addr[1] ), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15760_4_lut.init = 16'hc088;
    LUT4 i15759_4_lut (.A(div_factor_reg[25]), .B(\register_addr[1] ), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15759_4_lut.init = 16'hc088;
    LUT4 i15758_4_lut (.A(div_factor_reg[26]), .B(\register_addr[1] ), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n100[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15758_4_lut.init = 16'hc088;
    LUT4 i15757_4_lut (.A(div_factor_reg[27]), .B(\register_addr[1] ), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15757_4_lut.init = 16'hc088;
    LUT4 i15756_4_lut (.A(div_factor_reg[28]), .B(\register_addr[1] ), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15756_4_lut.init = 16'hc088;
    LUT4 i15755_4_lut (.A(div_factor_reg[29]), .B(\register_addr[1] ), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15755_4_lut.init = 16'hc088;
    LUT4 i15754_4_lut (.A(div_factor_reg[30]), .B(\register_addr[1] ), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15754_4_lut.init = 16'hc088;
    LUT4 i15753_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15753_4_lut.init = 16'hc088;
    LUT4 mux_1610_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n4121), 
         .Z(n4122[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n4121), .Z(n4122[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i7_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_329_4_lut (.A(rw), .B(n32181), .C(n32233), .D(n29750), 
         .Z(n32150)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i2_3_lut_rep_329_4_lut.init = 16'h0400;
    LUT4 mux_1610_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n4121), 
         .Z(n4122[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i20_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(rw), .B(n32181), .C(n32279), .D(n13118), 
         .Z(n4121)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i2_3_lut_4_lut.init = 16'h0400;
    LUT4 i23092_3_lut_3_lut_4_lut (.A(\register_addr[0] ), .B(n32231), .C(n32235), 
         .D(n32232), .Z(n22529)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(116[11:28])
    defparam i23092_3_lut_3_lut_4_lut.init = 16'h001f;
    LUT4 i8091_3_lut_4_lut_4_lut_4_lut (.A(\register_addr[0] ), .B(n32231), 
         .C(n32235), .D(n32232), .Z(n14812)) /* synthesis lut_function=(!(A (C+(D))+!A (B+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(116[11:28])
    defparam i8091_3_lut_4_lut_4_lut_4_lut.init = 16'h001b;
    LUT4 mux_1610_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n4121), .Z(n4122[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n4121), 
         .Z(n4122[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n4121), .Z(n4122[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i5_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 mux_1610_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n4121), .Z(n4122[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n4121), .Z(n4122[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n4121), 
         .Z(n4122[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n4121), .Z(n4122[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i2_3_lut.init = 16'hcaca;
    LUT4 i23134_2_lut_2_lut_3_lut_4_lut (.A(n32282), .B(\register_addr[1] ), 
         .C(n32314), .D(n32315), .Z(n30020)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i23134_2_lut_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i2_3_lut_4_lut_adj_26 (.A(n32282), .B(\register_addr[1] ), .C(n32305), 
         .D(n32315), .Z(n28426)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i2_3_lut_4_lut_adj_26.init = 16'h0040;
    LUT4 i23057_2_lut_2_lut_3_lut_4_lut (.A(n32282), .B(\register_addr[1] ), 
         .C(n32261), .D(n32315), .Z(n30019)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i23057_2_lut_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 equal_139_i15_2_lut_rep_366_3_lut_4_lut (.A(n32282), .B(\register_addr[1] ), 
         .C(n32232), .D(\register_addr[0] ), .Z(n32187)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam equal_139_i15_2_lut_rep_366_3_lut_4_lut.init = 16'hfffb;
    LUT4 mux_1610_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n4121), 
         .Z(n4122[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i17_3_lut.init = 16'hcaca;
    LUT4 i118_1_lut (.A(limit_c_0), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 mux_1610_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n4121), 
         .Z(n4122[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n4121), 
         .Z(n4122[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n4121), 
         .Z(n4122[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i14_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut (.A(n29750), .B(n32233), .C(n32159), .D(n34065), 
         .Z(n13444)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;
    defparam i1_2_lut_4_lut.init = 16'hff20;
    LUT4 mux_1610_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n4121), 
         .Z(n4122[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i25_3_lut.init = 16'hcaca;
    LUT4 i4412_3_lut (.A(prev_limit_latched), .B(n34065), .C(limit_latched), 
         .Z(n11127)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i4412_3_lut.init = 16'hdcdc;
    LUT4 mux_1610_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n4121), 
         .Z(n4122[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i28_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(n14419), .B(\register_addr[0] ), .C(n32232), .D(n32231), 
         .Z(n9478)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut.init = 16'h0008;
    LUT4 i15354_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n1_c)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15354_2_lut.init = 16'h2222;
    LUT4 mux_1918_Mux_3_i2_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), 
         .C(\register_addr[0] ), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1918_Mux_3_i2_3_lut.init = 16'hcaca;
    LUT4 i15353_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n1_adj_12)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15353_2_lut.init = 16'h2222;
    LUT4 mux_1918_Mux_4_i2_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), 
         .C(\register_addr[0] ), .Z(n2_adj_13)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1918_Mux_4_i2_3_lut.init = 16'hcaca;
    LUT4 i15352_2_lut (.A(Stepper_X_Dir_c), .B(\register_addr[0] ), .Z(n1_adj_14)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15352_2_lut.init = 16'h2222;
    LUT4 mux_1918_Mux_5_i2_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), 
         .C(\register_addr[0] ), .Z(n2_adj_15)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1918_Mux_5_i2_3_lut.init = 16'hcaca;
    LUT4 i15349_2_lut (.A(Stepper_X_En_c), .B(\register_addr[0] ), .Z(n1_adj_16)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15349_2_lut.init = 16'h2222;
    LUT4 mux_1918_Mux_6_i2_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), 
         .C(\register_addr[0] ), .Z(n2_adj_17)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1918_Mux_6_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1918_Mux_7_i2_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), 
         .C(\register_addr[0] ), .Z(n2_adj_18)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1918_Mux_7_i2_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n100[7]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n100[20]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n100[23]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n100[26]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    LUT4 i22866_3_lut (.A(Stepper_X_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n30369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22866_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n4121), 
         .Z(n4122[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i27_3_lut.init = 16'hcaca;
    LUT4 i22867_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n30370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22867_3_lut.init = 16'hcaca;
    PFUMX mux_1918_Mux_3_i3 (.BLUT(n1_c), .ALUT(n2), .C0(\register_addr[1] ), 
          .Z(n6439[3]));
    PFUMX mux_1918_Mux_4_i3 (.BLUT(n1_adj_12), .ALUT(n2_adj_13), .C0(\register_addr[1] ), 
          .Z(n100[4]));
    PFUMX mux_1918_Mux_5_i3 (.BLUT(n1_adj_14), .ALUT(n2_adj_15), .C0(\register_addr[1] ), 
          .Z(n100[5]));
    PFUMX mux_1918_Mux_6_i3 (.BLUT(n1_adj_16), .ALUT(n2_adj_17), .C0(\register_addr[1] ), 
          .Z(n100[6]));
    PFUMX mux_1918_Mux_7_i3 (.BLUT(n1), .ALUT(n2_adj_18), .C0(\register_addr[1] ), 
          .Z(n100[7]));
    PFUMX i22868 (.BLUT(n30369), .ALUT(n30370), .C0(\register_addr[1] ), 
          .Z(n30371));
    LUT4 i22896_3_lut (.A(Stepper_X_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n30399)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22896_3_lut.init = 16'hcaca;
    PFUMX i22898 (.BLUT(n30399), .ALUT(n30400), .C0(\register_addr[1] ), 
          .Z(n30401));
    LUT4 i22897_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n30400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22897_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i3 (.D(n6439[3]), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30395), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30401), .SP(n2769), .CD(n9485), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i22890_3_lut (.A(Stepper_X_M2_c_2), .B(n34), .C(\register_addr[0] ), 
         .Z(n30393)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22890_3_lut.init = 16'hcaca;
    LUT4 i22891_3_lut (.A(div_factor_reg[2]), .B(steps_reg[2]), .C(\register_addr[0] ), 
         .Z(n30394)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22891_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62_adj_21), .C(n58_adj_22), .D(n50_adj_23), 
         .Z(n28062)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[0]), .B(steps_reg[27]), .C(steps_reg[31]), 
         .D(steps_reg[30]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60_adj_24), .C(n54_adj_25), .D(n42_adj_26), 
         .Z(n62_adj_21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[15]), .B(n52_adj_27), .C(n38_adj_28), 
         .D(steps_reg[11]), .Z(n58_adj_22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[18]), .B(steps_reg[8]), .C(steps_reg[2]), 
         .D(steps_reg[16]), .Z(n50_adj_23)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[24]), .B(steps_reg[1]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[6]), .B(n56_adj_29), .C(n46_adj_30), 
         .D(steps_reg[10]), .Z(n60_adj_24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[7]), .B(steps_reg[26]), .C(steps_reg[25]), 
         .D(steps_reg[5]), .Z(n54_adj_25)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[4]), .B(steps_reg[21]), .Z(n42_adj_26)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[19]), .B(steps_reg[3]), .C(steps_reg[22]), 
         .D(steps_reg[13]), .Z(n56_adj_29)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[20]), .B(steps_reg[14]), .Z(n46_adj_30)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[29]), .B(steps_reg[12]), .C(steps_reg[9]), 
         .D(steps_reg[17]), .Z(n52_adj_27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[28]), .B(steps_reg[23]), .Z(n38_adj_28)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    IFS1P3DX fault_latched_178 (.D(Stepper_X_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1P3AX int_step_182 (.D(n32142), .SP(n24), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27430), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    LUT4 mux_1610_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n4121), 
         .Z(n4122[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i24_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27429), .COUT(n27430), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27428), .COUT(n27429), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27427), .COUT(n27428), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27426), .COUT(n27427), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    LUT4 mux_1610_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n4121), 
         .Z(n4122[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i32_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27425), .COUT(n27426), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27424), .COUT(n27425), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27423), .COUT(n27424), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    LUT4 mux_1610_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n4121), 
         .Z(n4122[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i31_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27422), .COUT(n27423), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27421), .COUT(n27422), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27420), .COUT(n27421), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27419), .COUT(n27420), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27418), .COUT(n27419), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27417), .COUT(n27418), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27416), .COUT(n27417), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27415), .COUT(n27416), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(step_clk), .C1(n34), .D1(prev_step_clk), 
          .COUT(n27415), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 mux_1610_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n4121), 
         .Z(n4122[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i30_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n13444), .CD(n34069), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=580, LSE_RLINE=593 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    LUT4 mux_1610_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n4121), 
         .Z(n4122[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n4121), 
         .Z(n4122[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n4121), 
         .Z(n4122[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1610_i22_3_lut.init = 16'hcaca;
    ClockDivider_U8 step_clk_gen (.GND_net(GND_net), .step_clk(step_clk), 
            .debug_c_c(debug_c_c), .n34066(n34066), .div_factor_reg({div_factor_reg}), 
            .n34065(n34065)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U8
//

module ClockDivider_U8 (GND_net, step_clk, debug_c_c, n34066, div_factor_reg, 
            n34065) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output step_clk;
    input debug_c_c;
    input n34066;
    input [31:0]div_factor_reg;
    input n34065;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n27648;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n27649, n27306;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n27307, n27305, n27647, n27304, n27303, n27302, n27301, 
        n27300, n27299, n27298, n7961, n27297, n27296, n27295, 
        n27294;
    wire [31:0]n40;
    
    wire n7996, n27494, n27493, n27293, n27492, n27491, n27490, 
        n27489, n27488, n27292, n27487, n27486, n27485, n27484, 
        n27291, n27483, n27482, n27481, n27290, n27480, n27479, 
        n27289, n32131, n27288, n27287, n27286, n27285, n27284, 
        n27283, n27282, n27281, n27280, n27279, n27278, n8030, 
        n27277, n27276, n16722, n27275, n27274, n27273, n27272, 
        n27271, n27270, n27269, n27268, n27267, n27266, n27265, 
        n27264, n27263, n27662, n27661, n27660, n27659, n27658, 
        n27310, n27657, n27656, n27655, n27654, n27309, n27653, 
        n27652, n27651, n27308, n27650;
    
    CCU2D count_2662_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27648), .COUT(n27649), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2662_add_4_5.INJECT1_0 = "NO";
    defparam count_2662_add_4_5.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27306), .COUT(n27307));
    defparam sub_2052_add_2_25.INIT0 = 16'h5999;
    defparam sub_2052_add_2_25.INIT1 = 16'h5999;
    defparam sub_2052_add_2_25.INJECT1_0 = "NO";
    defparam sub_2052_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27305), .COUT(n27306));
    defparam sub_2052_add_2_23.INIT0 = 16'h5999;
    defparam sub_2052_add_2_23.INIT1 = 16'h5999;
    defparam sub_2052_add_2_23.INJECT1_0 = "NO";
    defparam sub_2052_add_2_23.INJECT1_1 = "NO";
    CCU2D count_2662_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27647), .COUT(n27648), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2662_add_4_3.INJECT1_0 = "NO";
    defparam count_2662_add_4_3.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27304), .COUT(n27305));
    defparam sub_2052_add_2_21.INIT0 = 16'h5999;
    defparam sub_2052_add_2_21.INIT1 = 16'h5999;
    defparam sub_2052_add_2_21.INJECT1_0 = "NO";
    defparam sub_2052_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27303), .COUT(n27304));
    defparam sub_2052_add_2_19.INIT0 = 16'h5999;
    defparam sub_2052_add_2_19.INIT1 = 16'h5999;
    defparam sub_2052_add_2_19.INJECT1_0 = "NO";
    defparam sub_2052_add_2_19.INJECT1_1 = "NO";
    CCU2D count_2662_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27647), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_1.INIT0 = 16'hF000;
    defparam count_2662_add_4_1.INIT1 = 16'h0555;
    defparam count_2662_add_4_1.INJECT1_0 = "NO";
    defparam count_2662_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27302), .COUT(n27303));
    defparam sub_2052_add_2_17.INIT0 = 16'h5999;
    defparam sub_2052_add_2_17.INIT1 = 16'h5999;
    defparam sub_2052_add_2_17.INJECT1_0 = "NO";
    defparam sub_2052_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27301), .COUT(n27302));
    defparam sub_2052_add_2_15.INIT0 = 16'h5999;
    defparam sub_2052_add_2_15.INIT1 = 16'h5999;
    defparam sub_2052_add_2_15.INJECT1_0 = "NO";
    defparam sub_2052_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27300), .COUT(n27301));
    defparam sub_2052_add_2_13.INIT0 = 16'h5999;
    defparam sub_2052_add_2_13.INIT1 = 16'h5999;
    defparam sub_2052_add_2_13.INJECT1_0 = "NO";
    defparam sub_2052_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27299), .COUT(n27300));
    defparam sub_2052_add_2_11.INIT0 = 16'h5999;
    defparam sub_2052_add_2_11.INIT1 = 16'h5999;
    defparam sub_2052_add_2_11.INJECT1_0 = "NO";
    defparam sub_2052_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27298), .COUT(n27299));
    defparam sub_2052_add_2_9.INIT0 = 16'h5999;
    defparam sub_2052_add_2_9.INIT1 = 16'h5999;
    defparam sub_2052_add_2_9.INJECT1_0 = "NO";
    defparam sub_2052_add_2_9.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n7961), .CK(debug_c_c), .CD(n34066), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_2052_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27297), .COUT(n27298));
    defparam sub_2052_add_2_7.INIT0 = 16'h5999;
    defparam sub_2052_add_2_7.INIT1 = 16'h5999;
    defparam sub_2052_add_2_7.INJECT1_0 = "NO";
    defparam sub_2052_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27296), .COUT(n27297));
    defparam sub_2052_add_2_5.INIT0 = 16'h5999;
    defparam sub_2052_add_2_5.INIT1 = 16'h5999;
    defparam sub_2052_add_2_5.INJECT1_0 = "NO";
    defparam sub_2052_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27295), .COUT(n27296));
    defparam sub_2052_add_2_3.INIT0 = 16'h5999;
    defparam sub_2052_add_2_3.INIT1 = 16'h5999;
    defparam sub_2052_add_2_3.INJECT1_0 = "NO";
    defparam sub_2052_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27295));
    defparam sub_2052_add_2_1.INIT0 = 16'h0000;
    defparam sub_2052_add_2_1.INIT1 = 16'h5999;
    defparam sub_2052_add_2_1.INJECT1_0 = "NO";
    defparam sub_2052_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27294), .S1(n7996));
    defparam sub_2054_add_2_33.INIT0 = 16'h5999;
    defparam sub_2054_add_2_33.INIT1 = 16'h0000;
    defparam sub_2054_add_2_33.INJECT1_0 = "NO";
    defparam sub_2054_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27494), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27493), .COUT(n27494), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27293), .COUT(n27294));
    defparam sub_2054_add_2_31.INIT0 = 16'h5999;
    defparam sub_2054_add_2_31.INIT1 = 16'h5999;
    defparam sub_2054_add_2_31.INJECT1_0 = "NO";
    defparam sub_2054_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27492), .COUT(n27493), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27491), .COUT(n27492), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27490), .COUT(n27491), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27489), .COUT(n27490), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27488), .COUT(n27489), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27292), .COUT(n27293));
    defparam sub_2054_add_2_29.INIT0 = 16'h5999;
    defparam sub_2054_add_2_29.INIT1 = 16'h5999;
    defparam sub_2054_add_2_29.INJECT1_0 = "NO";
    defparam sub_2054_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27487), .COUT(n27488), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27486), .COUT(n27487), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27485), .COUT(n27486), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27484), .COUT(n27485), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27291), .COUT(n27292));
    defparam sub_2054_add_2_27.INIT0 = 16'h5999;
    defparam sub_2054_add_2_27.INIT1 = 16'h5999;
    defparam sub_2054_add_2_27.INJECT1_0 = "NO";
    defparam sub_2054_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27483), .COUT(n27484), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27482), .COUT(n27483), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27481), .COUT(n27482), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27290), .COUT(n27291));
    defparam sub_2054_add_2_25.INIT0 = 16'h5999;
    defparam sub_2054_add_2_25.INIT1 = 16'h5999;
    defparam sub_2054_add_2_25.INJECT1_0 = "NO";
    defparam sub_2054_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27480), .COUT(n27481), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27479), .COUT(n27480), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27289), .COUT(n27290));
    defparam sub_2054_add_2_23.INIT0 = 16'h5999;
    defparam sub_2054_add_2_23.INIT1 = 16'h5999;
    defparam sub_2054_add_2_23.INJECT1_0 = "NO";
    defparam sub_2054_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27479), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    FD1S3IX count_2662__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i0.GSR = "ENABLED";
    CCU2D sub_2054_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27288), .COUT(n27289));
    defparam sub_2054_add_2_21.INIT0 = 16'h5999;
    defparam sub_2054_add_2_21.INIT1 = 16'h5999;
    defparam sub_2054_add_2_21.INJECT1_0 = "NO";
    defparam sub_2054_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27287), .COUT(n27288));
    defparam sub_2054_add_2_19.INIT0 = 16'h5999;
    defparam sub_2054_add_2_19.INIT1 = 16'h5999;
    defparam sub_2054_add_2_19.INJECT1_0 = "NO";
    defparam sub_2054_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27286), .COUT(n27287));
    defparam sub_2054_add_2_17.INIT0 = 16'h5999;
    defparam sub_2054_add_2_17.INIT1 = 16'h5999;
    defparam sub_2054_add_2_17.INJECT1_0 = "NO";
    defparam sub_2054_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27285), .COUT(n27286));
    defparam sub_2054_add_2_15.INIT0 = 16'h5999;
    defparam sub_2054_add_2_15.INIT1 = 16'h5999;
    defparam sub_2054_add_2_15.INJECT1_0 = "NO";
    defparam sub_2054_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27284), .COUT(n27285));
    defparam sub_2054_add_2_13.INIT0 = 16'h5999;
    defparam sub_2054_add_2_13.INIT1 = 16'h5999;
    defparam sub_2054_add_2_13.INJECT1_0 = "NO";
    defparam sub_2054_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27283), .COUT(n27284));
    defparam sub_2054_add_2_11.INIT0 = 16'h5999;
    defparam sub_2054_add_2_11.INIT1 = 16'h5999;
    defparam sub_2054_add_2_11.INJECT1_0 = "NO";
    defparam sub_2054_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27282), .COUT(n27283));
    defparam sub_2054_add_2_9.INIT0 = 16'h5999;
    defparam sub_2054_add_2_9.INIT1 = 16'h5999;
    defparam sub_2054_add_2_9.INJECT1_0 = "NO";
    defparam sub_2054_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27281), .COUT(n27282));
    defparam sub_2054_add_2_7.INIT0 = 16'h5999;
    defparam sub_2054_add_2_7.INIT1 = 16'h5999;
    defparam sub_2054_add_2_7.INJECT1_0 = "NO";
    defparam sub_2054_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27280), .COUT(n27281));
    defparam sub_2054_add_2_5.INIT0 = 16'h5999;
    defparam sub_2054_add_2_5.INIT1 = 16'h5999;
    defparam sub_2054_add_2_5.INJECT1_0 = "NO";
    defparam sub_2054_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27279), .COUT(n27280));
    defparam sub_2054_add_2_3.INIT0 = 16'h5999;
    defparam sub_2054_add_2_3.INIT1 = 16'h5999;
    defparam sub_2054_add_2_3.INJECT1_0 = "NO";
    defparam sub_2054_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2054_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27279));
    defparam sub_2054_add_2_1.INIT0 = 16'h0000;
    defparam sub_2054_add_2_1.INIT1 = 16'h5999;
    defparam sub_2054_add_2_1.INJECT1_0 = "NO";
    defparam sub_2054_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27278), .S1(n8030));
    defparam sub_2055_add_2_33.INIT0 = 16'hf555;
    defparam sub_2055_add_2_33.INIT1 = 16'h0000;
    defparam sub_2055_add_2_33.INJECT1_0 = "NO";
    defparam sub_2055_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27277), .COUT(n27278));
    defparam sub_2055_add_2_31.INIT0 = 16'hf555;
    defparam sub_2055_add_2_31.INIT1 = 16'hf555;
    defparam sub_2055_add_2_31.INJECT1_0 = "NO";
    defparam sub_2055_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27276), .COUT(n27277));
    defparam sub_2055_add_2_29.INIT0 = 16'hf555;
    defparam sub_2055_add_2_29.INIT1 = 16'hf555;
    defparam sub_2055_add_2_29.INJECT1_0 = "NO";
    defparam sub_2055_add_2_29.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n32131), .PD(n16722), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_2055_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27275), .COUT(n27276));
    defparam sub_2055_add_2_27.INIT0 = 16'hf555;
    defparam sub_2055_add_2_27.INIT1 = 16'hf555;
    defparam sub_2055_add_2_27.INJECT1_0 = "NO";
    defparam sub_2055_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27274), .COUT(n27275));
    defparam sub_2055_add_2_25.INIT0 = 16'hf555;
    defparam sub_2055_add_2_25.INIT1 = 16'hf555;
    defparam sub_2055_add_2_25.INJECT1_0 = "NO";
    defparam sub_2055_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27273), .COUT(n27274));
    defparam sub_2055_add_2_23.INIT0 = 16'hf555;
    defparam sub_2055_add_2_23.INIT1 = 16'hf555;
    defparam sub_2055_add_2_23.INJECT1_0 = "NO";
    defparam sub_2055_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27272), .COUT(n27273));
    defparam sub_2055_add_2_21.INIT0 = 16'hf555;
    defparam sub_2055_add_2_21.INIT1 = 16'hf555;
    defparam sub_2055_add_2_21.INJECT1_0 = "NO";
    defparam sub_2055_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27271), .COUT(n27272));
    defparam sub_2055_add_2_19.INIT0 = 16'hf555;
    defparam sub_2055_add_2_19.INIT1 = 16'hf555;
    defparam sub_2055_add_2_19.INJECT1_0 = "NO";
    defparam sub_2055_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27270), .COUT(n27271));
    defparam sub_2055_add_2_17.INIT0 = 16'hf555;
    defparam sub_2055_add_2_17.INIT1 = 16'hf555;
    defparam sub_2055_add_2_17.INJECT1_0 = "NO";
    defparam sub_2055_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27269), .COUT(n27270));
    defparam sub_2055_add_2_15.INIT0 = 16'hf555;
    defparam sub_2055_add_2_15.INIT1 = 16'hf555;
    defparam sub_2055_add_2_15.INJECT1_0 = "NO";
    defparam sub_2055_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27268), .COUT(n27269));
    defparam sub_2055_add_2_13.INIT0 = 16'hf555;
    defparam sub_2055_add_2_13.INIT1 = 16'hf555;
    defparam sub_2055_add_2_13.INJECT1_0 = "NO";
    defparam sub_2055_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27267), .COUT(n27268));
    defparam sub_2055_add_2_11.INIT0 = 16'hf555;
    defparam sub_2055_add_2_11.INIT1 = 16'hf555;
    defparam sub_2055_add_2_11.INJECT1_0 = "NO";
    defparam sub_2055_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27266), .COUT(n27267));
    defparam sub_2055_add_2_9.INIT0 = 16'hf555;
    defparam sub_2055_add_2_9.INIT1 = 16'hf555;
    defparam sub_2055_add_2_9.INJECT1_0 = "NO";
    defparam sub_2055_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27265), .COUT(n27266));
    defparam sub_2055_add_2_7.INIT0 = 16'hf555;
    defparam sub_2055_add_2_7.INIT1 = 16'hf555;
    defparam sub_2055_add_2_7.INJECT1_0 = "NO";
    defparam sub_2055_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27264), .COUT(n27265));
    defparam sub_2055_add_2_5.INIT0 = 16'hf555;
    defparam sub_2055_add_2_5.INIT1 = 16'hf555;
    defparam sub_2055_add_2_5.INJECT1_0 = "NO";
    defparam sub_2055_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27263), .COUT(n27264));
    defparam sub_2055_add_2_3.INIT0 = 16'hf555;
    defparam sub_2055_add_2_3.INIT1 = 16'hf555;
    defparam sub_2055_add_2_3.INJECT1_0 = "NO";
    defparam sub_2055_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2055_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27263));
    defparam sub_2055_add_2_1.INIT0 = 16'h0000;
    defparam sub_2055_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2055_add_2_1.INJECT1_0 = "NO";
    defparam sub_2055_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n32131), .CD(n16722), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    FD1S3IX count_2662__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i1.GSR = "ENABLED";
    FD1S3IX count_2662__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i2.GSR = "ENABLED";
    FD1S3IX count_2662__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i3.GSR = "ENABLED";
    FD1S3IX count_2662__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i4.GSR = "ENABLED";
    FD1S3IX count_2662__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i5.GSR = "ENABLED";
    FD1S3IX count_2662__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i6.GSR = "ENABLED";
    FD1S3IX count_2662__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i7.GSR = "ENABLED";
    FD1S3IX count_2662__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i8.GSR = "ENABLED";
    FD1S3IX count_2662__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i9.GSR = "ENABLED";
    FD1S3IX count_2662__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i10.GSR = "ENABLED";
    FD1S3IX count_2662__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i11.GSR = "ENABLED";
    FD1S3IX count_2662__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i12.GSR = "ENABLED";
    FD1S3IX count_2662__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i13.GSR = "ENABLED";
    FD1S3IX count_2662__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i14.GSR = "ENABLED";
    FD1S3IX count_2662__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i15.GSR = "ENABLED";
    FD1S3IX count_2662__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i16.GSR = "ENABLED";
    FD1S3IX count_2662__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i17.GSR = "ENABLED";
    FD1S3IX count_2662__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i18.GSR = "ENABLED";
    FD1S3IX count_2662__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i19.GSR = "ENABLED";
    FD1S3IX count_2662__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i20.GSR = "ENABLED";
    FD1S3IX count_2662__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i21.GSR = "ENABLED";
    FD1S3IX count_2662__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i22.GSR = "ENABLED";
    FD1S3IX count_2662__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i23.GSR = "ENABLED";
    FD1S3IX count_2662__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i24.GSR = "ENABLED";
    FD1S3IX count_2662__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i25.GSR = "ENABLED";
    FD1S3IX count_2662__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i26.GSR = "ENABLED";
    FD1S3IX count_2662__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i27.GSR = "ENABLED";
    FD1S3IX count_2662__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i28.GSR = "ENABLED";
    FD1S3IX count_2662__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i29.GSR = "ENABLED";
    FD1S3IX count_2662__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i30.GSR = "ENABLED";
    FD1S3IX count_2662__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n32131), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662__i31.GSR = "ENABLED";
    LUT4 i1020_2_lut_rep_310 (.A(n7996), .B(n34065), .Z(n32131)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i1020_2_lut_rep_310.init = 16'heeee;
    LUT4 i10030_2_lut_3_lut (.A(n7996), .B(n34065), .C(n8030), .Z(n16722)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i10030_2_lut_3_lut.init = 16'he0e0;
    CCU2D count_2662_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27662), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_33.INIT1 = 16'h0000;
    defparam count_2662_add_4_33.INJECT1_0 = "NO";
    defparam count_2662_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2662_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27661), .COUT(n27662), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2662_add_4_31.INJECT1_0 = "NO";
    defparam count_2662_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2662_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27660), .COUT(n27661), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2662_add_4_29.INJECT1_0 = "NO";
    defparam count_2662_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2662_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27659), .COUT(n27660), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2662_add_4_27.INJECT1_0 = "NO";
    defparam count_2662_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2662_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27658), .COUT(n27659), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2662_add_4_25.INJECT1_0 = "NO";
    defparam count_2662_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27310), .S1(n7961));
    defparam sub_2052_add_2_33.INIT0 = 16'h5555;
    defparam sub_2052_add_2_33.INIT1 = 16'h0000;
    defparam sub_2052_add_2_33.INJECT1_0 = "NO";
    defparam sub_2052_add_2_33.INJECT1_1 = "NO";
    CCU2D count_2662_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27657), .COUT(n27658), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2662_add_4_23.INJECT1_0 = "NO";
    defparam count_2662_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2662_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27656), .COUT(n27657), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2662_add_4_21.INJECT1_0 = "NO";
    defparam count_2662_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2662_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27655), .COUT(n27656), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2662_add_4_19.INJECT1_0 = "NO";
    defparam count_2662_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2662_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27654), .COUT(n27655), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2662_add_4_17.INJECT1_0 = "NO";
    defparam count_2662_add_4_17.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27309), .COUT(n27310));
    defparam sub_2052_add_2_31.INIT0 = 16'h5999;
    defparam sub_2052_add_2_31.INIT1 = 16'h5999;
    defparam sub_2052_add_2_31.INJECT1_0 = "NO";
    defparam sub_2052_add_2_31.INJECT1_1 = "NO";
    CCU2D count_2662_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27653), .COUT(n27654), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2662_add_4_15.INJECT1_0 = "NO";
    defparam count_2662_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2662_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27652), .COUT(n27653), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2662_add_4_13.INJECT1_0 = "NO";
    defparam count_2662_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2662_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27651), .COUT(n27652), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2662_add_4_11.INJECT1_0 = "NO";
    defparam count_2662_add_4_11.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27308), .COUT(n27309));
    defparam sub_2052_add_2_29.INIT0 = 16'h5999;
    defparam sub_2052_add_2_29.INIT1 = 16'h5999;
    defparam sub_2052_add_2_29.INJECT1_0 = "NO";
    defparam sub_2052_add_2_29.INJECT1_1 = "NO";
    CCU2D count_2662_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27650), .COUT(n27651), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2662_add_4_9.INJECT1_0 = "NO";
    defparam count_2662_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2662_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27649), .COUT(n27650), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2662_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2662_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2662_add_4_7.INJECT1_0 = "NO";
    defparam count_2662_add_4_7.INJECT1_1 = "NO";
    CCU2D sub_2052_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27307), .COUT(n27308));
    defparam sub_2052_add_2_27.INIT0 = 16'h5999;
    defparam sub_2052_add_2_27.INIT1 = 16'h5999;
    defparam sub_2052_add_2_27.INJECT1_0 = "NO";
    defparam sub_2052_add_2_27.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module EncoderPeripheral
//

module EncoderPeripheral (\read_size[0] , debug_c_c, n178, n32157, n32202, 
            read_value, prev_select, n32178, \register_addr[0] , n32235, 
            n32232, prev_select_adj_8, n30270, n32315, n29983, n32138, 
            n29977, n9, \read_size[2] , \register_addr[1] , n32282, 
            n32166, n32279, n32204, n32181, rw, n32149, n34065, 
            n32159, n13511, encoder_ra_c, encoder_rb_c, encoder_ri_c, 
            n14493, n14419, n32231, n16516, n16515, n6, n13588, 
            qreset, VCC_net, GND_net, \quadB_delayed[1] , \quadA_delayed[1] ) /* synthesis syn_module_defined=1 */ ;
    output \read_size[0] ;
    input debug_c_c;
    input n178;
    input n32157;
    input n32202;
    output [31:0]read_value;
    output prev_select;
    input n32178;
    input \register_addr[0] ;
    input n32235;
    input n32232;
    input prev_select_adj_8;
    output n30270;
    input n32315;
    input n29983;
    output n32138;
    input n29977;
    output n9;
    output \read_size[2] ;
    input \register_addr[1] ;
    input n32282;
    output n32166;
    input n32279;
    output n32204;
    input n32181;
    input rw;
    output n32149;
    input n34065;
    input n32159;
    output n13511;
    input encoder_ra_c;
    input encoder_rb_c;
    input encoder_ri_c;
    output n14493;
    input n14419;
    input n32231;
    output n16516;
    output n16515;
    output n6;
    input n13588;
    input qreset;
    input VCC_net;
    input GND_net;
    output \quadB_delayed[1] ;
    output \quadA_delayed[1] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [31:0]n100;
    wire [1:0]n1;
    wire [31:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(58[14:22])
    
    FD1P3IX read_size__i1 (.D(n32202), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n100[0]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1S3AX prev_select_126 (.D(n32178), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam prev_select_126.GSR = "ENABLED";
    FD1P3IX read_value__i31 (.D(n100[31]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_value__i30 (.D(n100[30]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n100[29]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n100[28]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n100[27]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n100[26]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n100[25]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n100[24]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n100[23]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n100[22]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n100[21]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n100[20]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n100[19]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n100[16]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n100[14]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n100[13]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n100[12]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n100[11]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n100[10]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n100[9]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n100[8]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n100[7]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n100[6]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n100[5]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n100[4]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n100[3]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n100[2]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n100[1]), .SP(n178), .CD(n32157), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i22767_2_lut_3_lut_3_lut_4_lut (.A(\register_addr[0] ), .B(n32235), 
         .C(n32232), .D(prev_select_adj_8), .Z(n30270)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[21:41])
    defparam i22767_2_lut_3_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_317_3_lut_3_lut_4_lut (.A(\register_addr[0] ), .B(n32235), 
         .C(n32315), .D(n29983), .Z(n32138)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[21:41])
    defparam i1_2_lut_rep_317_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i3_2_lut_3_lut_3_lut_4_lut (.A(\register_addr[0] ), .B(n32235), 
         .C(n32315), .D(n29977), .Z(n9)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[21:41])
    defparam i3_2_lut_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i15664_2_lut_4_lut_4_lut_4_lut (.A(\register_addr[0] ), .B(n32235), 
         .C(prev_select), .D(n32178), .Z(n1[1])) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[21:41])
    defparam i15664_2_lut_4_lut_4_lut_4_lut.init = 16'he2ee;
    FD1P3AX read_size__i2 (.D(n1[1]), .SP(n178), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=20, LSE_RCOL=47, LSE_LLINE=682, LSE_RLINE=692 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(72[9] 88[6])
    defparam read_size__i2.GSR = "ENABLED";
    LUT4 i2_2_lut_rep_345_2_lut_3_lut_4_lut (.A(\register_addr[1] ), .B(n32282), 
         .C(n32315), .D(\register_addr[0] ), .Z(n32166)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(77[9:33])
    defparam i2_2_lut_rep_345_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_383_3_lut_4_lut (.A(\register_addr[1] ), .B(n32282), 
         .C(n32279), .D(n32315), .Z(n32204)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(77[9:33])
    defparam i1_2_lut_rep_383_3_lut_4_lut.init = 16'hfffe;
    LUT4 i15022_2_lut (.A(\register[1] [0]), .B(\register_addr[0] ), .Z(n100[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15022_2_lut.init = 16'h8888;
    LUT4 i23095_3_lut_rep_328_4_lut_4_lut (.A(n32202), .B(n32232), .C(n32181), 
         .D(rw), .Z(n32149)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[21:41])
    defparam i23095_3_lut_rep_328_4_lut_4_lut.init = 16'h0020;
    LUT4 i23097_2_lut_4_lut_4_lut (.A(n32202), .B(n34065), .C(n32232), 
         .D(n32159), .Z(n13511)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[21:41])
    defparam i23097_2_lut_4_lut_4_lut.init = 16'hcecc;
    LUT4 i15192_2_lut (.A(\register[1] [31]), .B(\register_addr[0] ), .Z(n100[31])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15192_2_lut.init = 16'h8888;
    LUT4 i15194_2_lut (.A(\register[1] [30]), .B(\register_addr[0] ), .Z(n100[30])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15194_2_lut.init = 16'h8888;
    LUT4 i15196_2_lut (.A(\register[1] [29]), .B(\register_addr[0] ), .Z(n100[29])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15196_2_lut.init = 16'h8888;
    LUT4 i15197_2_lut (.A(\register[1] [28]), .B(\register_addr[0] ), .Z(n100[28])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15197_2_lut.init = 16'h8888;
    LUT4 i15198_2_lut (.A(\register[1] [27]), .B(\register_addr[0] ), .Z(n100[27])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15198_2_lut.init = 16'h8888;
    LUT4 i15199_2_lut (.A(\register[1] [26]), .B(\register_addr[0] ), .Z(n100[26])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15199_2_lut.init = 16'h8888;
    LUT4 i15200_2_lut (.A(\register[1] [25]), .B(\register_addr[0] ), .Z(n100[25])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15200_2_lut.init = 16'h8888;
    LUT4 i15201_2_lut (.A(\register[1] [24]), .B(\register_addr[0] ), .Z(n100[24])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15201_2_lut.init = 16'h8888;
    LUT4 i15206_2_lut (.A(\register[1] [23]), .B(\register_addr[0] ), .Z(n100[23])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15206_2_lut.init = 16'h8888;
    LUT4 i15209_2_lut (.A(\register[1] [22]), .B(\register_addr[0] ), .Z(n100[22])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15209_2_lut.init = 16'h8888;
    LUT4 i15210_2_lut (.A(\register[1] [21]), .B(\register_addr[0] ), .Z(n100[21])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15210_2_lut.init = 16'h8888;
    LUT4 i15211_2_lut (.A(\register[1] [20]), .B(\register_addr[0] ), .Z(n100[20])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15211_2_lut.init = 16'h8888;
    LUT4 i15212_2_lut (.A(\register[1] [19]), .B(\register_addr[0] ), .Z(n100[19])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15212_2_lut.init = 16'h8888;
    LUT4 i15213_2_lut (.A(\register[1] [18]), .B(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15213_2_lut.init = 16'h8888;
    LUT4 i15214_2_lut (.A(\register[1] [17]), .B(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15214_2_lut.init = 16'h8888;
    LUT4 i15215_2_lut (.A(\register[1] [16]), .B(\register_addr[0] ), .Z(n100[16])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15215_2_lut.init = 16'h8888;
    LUT4 i15216_2_lut (.A(\register[1] [15]), .B(\register_addr[0] ), .Z(n100[15])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15216_2_lut.init = 16'h8888;
    LUT4 i15217_2_lut (.A(\register[1] [14]), .B(\register_addr[0] ), .Z(n100[14])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15217_2_lut.init = 16'h8888;
    LUT4 i15218_2_lut (.A(\register[1] [13]), .B(\register_addr[0] ), .Z(n100[13])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15218_2_lut.init = 16'h8888;
    LUT4 i15219_2_lut (.A(\register[1] [12]), .B(\register_addr[0] ), .Z(n100[12])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15219_2_lut.init = 16'h8888;
    LUT4 i15220_2_lut (.A(\register[1] [11]), .B(\register_addr[0] ), .Z(n100[11])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15220_2_lut.init = 16'h8888;
    LUT4 i15221_2_lut (.A(\register[1] [10]), .B(\register_addr[0] ), .Z(n100[10])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15221_2_lut.init = 16'h8888;
    LUT4 i15223_2_lut (.A(\register[1] [9]), .B(\register_addr[0] ), .Z(n100[9])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15223_2_lut.init = 16'h8888;
    LUT4 i15224_2_lut (.A(\register[1] [8]), .B(\register_addr[0] ), .Z(n100[8])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15224_2_lut.init = 16'h8888;
    LUT4 i15227_2_lut (.A(\register[1] [7]), .B(\register_addr[0] ), .Z(n100[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15227_2_lut.init = 16'h8888;
    LUT4 i15228_2_lut (.A(\register[1] [6]), .B(\register_addr[0] ), .Z(n100[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15228_2_lut.init = 16'h8888;
    LUT4 i15229_2_lut (.A(\register[1] [5]), .B(\register_addr[0] ), .Z(n100[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15229_2_lut.init = 16'h8888;
    LUT4 i15230_2_lut (.A(\register[1] [4]), .B(\register_addr[0] ), .Z(n100[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam i15230_2_lut.init = 16'h8888;
    LUT4 mux_115_Mux_3_i1_3_lut (.A(encoder_ra_c), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n100[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_2_i1_3_lut (.A(encoder_rb_c), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n100[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_115_Mux_1_i1_3_lut (.A(encoder_ri_c), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n100[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(79[31:44])
    defparam mux_115_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n32202), .B(n29983), .C(n34065), 
         .D(n32315), .Z(n14493)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[21:41])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hf0f8;
    LUT4 i9795_2_lut_4_lut_4_lut (.A(n32202), .B(n14419), .C(n32231), 
         .D(n32232), .Z(n16516)) /* synthesis lut_function=(!(A ((D)+!B)+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[21:41])
    defparam i9795_2_lut_4_lut_4_lut.init = 16'h008c;
    LUT4 i9794_2_lut_4_lut_4_lut (.A(n32202), .B(n14419), .C(n32231), 
         .D(n32232), .Z(n16515)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(80[21:41])
    defparam i9794_2_lut_4_lut_4_lut.init = 16'hcc40;
    QuadratureDecoder q (.n6(n6), .debug_c_c(debug_c_c), .n13588(n13588), 
            .qreset(qreset), .\register[1] ({\register[1] }), .VCC_net(VCC_net), 
            .GND_net(GND_net), .encoder_rb_c(encoder_rb_c), .encoder_ra_c(encoder_ra_c), 
            .\quadB_delayed[1] (\quadB_delayed[1] ), .\quadA_delayed[1] (\quadA_delayed[1] )) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(92[20] 96[37])
    
endmodule
//
// Verilog Description of module QuadratureDecoder
//

module QuadratureDecoder (n6, debug_c_c, n13588, qreset, \register[1] , 
            VCC_net, GND_net, encoder_rb_c, encoder_ra_c, \quadB_delayed[1] , 
            \quadA_delayed[1] ) /* synthesis syn_module_defined=1 */ ;
    output n6;
    input debug_c_c;
    input n13588;
    input qreset;
    output [31:0]\register[1] ;
    input VCC_net;
    input GND_net;
    input encoder_rb_c;
    input encoder_ra_c;
    output \quadB_delayed[1] ;
    output \quadA_delayed[1] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    wire [2:0]quadB_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[27:40])
    wire [2:0]quadA_delayed;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(16[12:25])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(15[13:18])
    wire [31:0]n100;
    
    wire n27133, n27132, n27131, n27130, n27129, n27128, n27127, 
        n27126, n27125, n27124, n27123, n27122, n27121, n27120, 
        n27119, n27118;
    
    LUT4 i2_2_lut (.A(quadB_delayed[2]), .B(quadA_delayed[2]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(18[22:95])
    defparam i2_2_lut.init = 16'h6666;
    FD1P3IX count__i0 (.D(n100[0]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i0.GSR = "ENABLED";
    FD1P3IX count__i31 (.D(n100[31]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i31.GSR = "ENABLED";
    FD1P3IX count__i30 (.D(n100[30]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i30.GSR = "ENABLED";
    FD1P3IX count__i29 (.D(n100[29]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i29.GSR = "ENABLED";
    FD1P3IX count__i28 (.D(n100[28]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i28.GSR = "ENABLED";
    FD1P3IX count__i27 (.D(n100[27]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i27.GSR = "ENABLED";
    FD1P3IX count__i26 (.D(n100[26]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i26.GSR = "ENABLED";
    FD1P3IX count__i25 (.D(n100[25]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i25.GSR = "ENABLED";
    FD1P3IX count__i24 (.D(n100[24]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i24.GSR = "ENABLED";
    FD1P3IX count__i23 (.D(n100[23]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i23.GSR = "ENABLED";
    FD1P3IX count__i22 (.D(n100[22]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i22.GSR = "ENABLED";
    FD1P3IX count__i21 (.D(n100[21]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i21.GSR = "ENABLED";
    FD1P3IX count__i20 (.D(n100[20]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i20.GSR = "ENABLED";
    FD1P3IX count__i19 (.D(n100[19]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i19.GSR = "ENABLED";
    FD1P3IX count__i18 (.D(n100[18]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i18.GSR = "ENABLED";
    FD1P3IX count__i17 (.D(n100[17]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i17.GSR = "ENABLED";
    FD1P3IX count__i16 (.D(n100[16]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i16.GSR = "ENABLED";
    FD1P3IX count__i15 (.D(n100[15]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i15.GSR = "ENABLED";
    FD1P3IX count__i14 (.D(n100[14]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i14.GSR = "ENABLED";
    FD1P3IX count__i13 (.D(n100[13]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i13.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n100[12]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i12.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n100[11]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n100[10]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n100[9]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n100[8]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n100[7]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n100[6]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n100[5]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n100[4]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n100[3]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n100[2]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n100[1]), .SP(n13588), .CD(qreset), .CK(debug_c_c), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count__i1.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i0 (.D(count[0]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i0.GSR = "ENABLED";
    IFS1P3DX quadB_delayed_i0 (.D(encoder_rb_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadB_delayed[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i0.GSR = "ENABLED";
    IFS1P3DX quadA_delayed_i0 (.D(encoder_ra_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(quadA_delayed[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i0.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i1 (.D(count[1]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i1.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i2 (.D(count[2]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i2.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i3 (.D(count[3]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i3.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i4 (.D(count[4]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i4.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i5 (.D(count[5]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i5.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i6 (.D(count[6]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i6.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i7 (.D(count[7]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i7.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i8 (.D(count[8]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i8.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i9 (.D(count[9]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i9.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i10 (.D(count[10]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i10.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i11 (.D(count[11]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i11.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i12 (.D(count[12]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i12.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i13 (.D(count[13]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i13.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i14 (.D(count[14]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i14.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i15 (.D(count[15]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i15.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i16 (.D(count[16]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i16.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i17 (.D(count[17]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i17.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i18 (.D(count[18]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i18.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i19 (.D(count[19]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i19.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i20 (.D(count[20]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i20.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i21 (.D(count[21]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i21.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i22 (.D(count[22]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i22.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i23 (.D(count[23]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i23.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i24 (.D(count[24]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i24.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i25 (.D(count[25]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i25.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i26 (.D(count[26]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i26.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i27 (.D(count[27]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i27.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i28 (.D(count[28]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i28.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i29 (.D(count[29]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i29.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i30 (.D(count[30]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i30.GSR = "ENABLED";
    FD1P3AX count_at_reset_i0_i31 (.D(count[31]), .SP(qreset), .CK(debug_c_c), 
            .Q(\register[1] [31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam count_at_reset_i0_i31.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i1 (.D(quadB_delayed[0]), .CK(debug_c_c), .Q(\quadB_delayed[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadB_delayed_i2 (.D(\quadB_delayed[1] ), .CK(debug_c_c), .Q(quadB_delayed[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadB_delayed_i2.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i1 (.D(quadA_delayed[0]), .CK(debug_c_c), .Q(\quadA_delayed[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i1.GSR = "ENABLED";
    FD1S3AX quadA_delayed_i2 (.D(\quadA_delayed[1] ), .CK(debug_c_c), .Q(quadA_delayed[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=20, LSE_RCOL=37, LSE_LLINE=92, LSE_RLINE=96 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(21[9] 37[6])
    defparam quadA_delayed_i2.GSR = "ENABLED";
    CCU2D add_1706_33 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[30]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[31]), .D1(GND_net), .CIN(n27133), .S0(n100[30]), 
          .S1(n100[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_33.INIT0 = 16'h6969;
    defparam add_1706_33.INIT1 = 16'h6969;
    defparam add_1706_33.INJECT1_0 = "NO";
    defparam add_1706_33.INJECT1_1 = "NO";
    CCU2D add_1706_31 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[28]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[29]), .D1(GND_net), .CIN(n27132), .COUT(n27133), 
          .S0(n100[28]), .S1(n100[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_31.INIT0 = 16'h6969;
    defparam add_1706_31.INIT1 = 16'h6969;
    defparam add_1706_31.INJECT1_0 = "NO";
    defparam add_1706_31.INJECT1_1 = "NO";
    CCU2D add_1706_29 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[26]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[27]), .D1(GND_net), .CIN(n27131), .COUT(n27132), 
          .S0(n100[26]), .S1(n100[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_29.INIT0 = 16'h6969;
    defparam add_1706_29.INIT1 = 16'h6969;
    defparam add_1706_29.INJECT1_0 = "NO";
    defparam add_1706_29.INJECT1_1 = "NO";
    CCU2D add_1706_27 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[24]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[25]), .D1(GND_net), .CIN(n27130), .COUT(n27131), 
          .S0(n100[24]), .S1(n100[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_27.INIT0 = 16'h6969;
    defparam add_1706_27.INIT1 = 16'h6969;
    defparam add_1706_27.INJECT1_0 = "NO";
    defparam add_1706_27.INJECT1_1 = "NO";
    CCU2D add_1706_25 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[22]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[23]), .D1(GND_net), .CIN(n27129), .COUT(n27130), 
          .S0(n100[22]), .S1(n100[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_25.INIT0 = 16'h6969;
    defparam add_1706_25.INIT1 = 16'h6969;
    defparam add_1706_25.INJECT1_0 = "NO";
    defparam add_1706_25.INJECT1_1 = "NO";
    CCU2D add_1706_23 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[20]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[21]), .D1(GND_net), .CIN(n27128), .COUT(n27129), 
          .S0(n100[20]), .S1(n100[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_23.INIT0 = 16'h6969;
    defparam add_1706_23.INIT1 = 16'h6969;
    defparam add_1706_23.INJECT1_0 = "NO";
    defparam add_1706_23.INJECT1_1 = "NO";
    CCU2D add_1706_21 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[18]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[19]), .D1(GND_net), .CIN(n27127), .COUT(n27128), 
          .S0(n100[18]), .S1(n100[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_21.INIT0 = 16'h6969;
    defparam add_1706_21.INIT1 = 16'h6969;
    defparam add_1706_21.INJECT1_0 = "NO";
    defparam add_1706_21.INJECT1_1 = "NO";
    CCU2D add_1706_19 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[16]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[17]), .D1(GND_net), .CIN(n27126), .COUT(n27127), 
          .S0(n100[16]), .S1(n100[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_19.INIT0 = 16'h6969;
    defparam add_1706_19.INIT1 = 16'h6969;
    defparam add_1706_19.INJECT1_0 = "NO";
    defparam add_1706_19.INJECT1_1 = "NO";
    CCU2D add_1706_17 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[14]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[15]), .D1(GND_net), .CIN(n27125), .COUT(n27126), 
          .S0(n100[14]), .S1(n100[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_17.INIT0 = 16'h6969;
    defparam add_1706_17.INIT1 = 16'h6969;
    defparam add_1706_17.INJECT1_0 = "NO";
    defparam add_1706_17.INJECT1_1 = "NO";
    CCU2D add_1706_15 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[12]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[13]), .D1(GND_net), .CIN(n27124), .COUT(n27125), 
          .S0(n100[12]), .S1(n100[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_15.INIT0 = 16'h6969;
    defparam add_1706_15.INIT1 = 16'h6969;
    defparam add_1706_15.INJECT1_0 = "NO";
    defparam add_1706_15.INJECT1_1 = "NO";
    CCU2D add_1706_13 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[10]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[11]), .D1(GND_net), .CIN(n27123), .COUT(n27124), 
          .S0(n100[10]), .S1(n100[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_13.INIT0 = 16'h6969;
    defparam add_1706_13.INIT1 = 16'h6969;
    defparam add_1706_13.INJECT1_0 = "NO";
    defparam add_1706_13.INJECT1_1 = "NO";
    CCU2D add_1706_11 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[8]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[9]), .D1(GND_net), .CIN(n27122), .COUT(n27123), 
          .S0(n100[8]), .S1(n100[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_11.INIT0 = 16'h6969;
    defparam add_1706_11.INIT1 = 16'h6969;
    defparam add_1706_11.INJECT1_0 = "NO";
    defparam add_1706_11.INJECT1_1 = "NO";
    CCU2D add_1706_9 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[6]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[7]), .D1(GND_net), .CIN(n27121), .COUT(n27122), 
          .S0(n100[6]), .S1(n100[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_9.INIT0 = 16'h6969;
    defparam add_1706_9.INIT1 = 16'h6969;
    defparam add_1706_9.INJECT1_0 = "NO";
    defparam add_1706_9.INJECT1_1 = "NO";
    CCU2D add_1706_7 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[4]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[5]), .D1(GND_net), .CIN(n27120), .COUT(n27121), 
          .S0(n100[4]), .S1(n100[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_7.INIT0 = 16'h6969;
    defparam add_1706_7.INIT1 = 16'h6969;
    defparam add_1706_7.INJECT1_0 = "NO";
    defparam add_1706_7.INJECT1_1 = "NO";
    CCU2D add_1706_5 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[2]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[3]), .D1(GND_net), .CIN(n27119), .COUT(n27120), 
          .S0(n100[2]), .S1(n100[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_5.INIT0 = 16'h6969;
    defparam add_1706_5.INIT1 = 16'h6969;
    defparam add_1706_5.INJECT1_0 = "NO";
    defparam add_1706_5.INJECT1_1 = "NO";
    CCU2D add_1706_3 (.A0(\quadA_delayed[1] ), .B0(quadB_delayed[2]), .C0(count[0]), 
          .D0(GND_net), .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), 
          .C1(count[1]), .D1(GND_net), .CIN(n27118), .COUT(n27119), 
          .S0(n100[0]), .S1(n100[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_3.INIT0 = 16'h9696;
    defparam add_1706_3.INIT1 = 16'h6969;
    defparam add_1706_3.INJECT1_0 = "NO";
    defparam add_1706_3.INJECT1_1 = "NO";
    CCU2D add_1706_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\quadA_delayed[1] ), .B1(quadB_delayed[2]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27118));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/encoder.v(31[5] 36[8])
    defparam add_1706_1.INIT0 = 16'hF000;
    defparam add_1706_1.INIT1 = 16'h6666;
    defparam add_1706_1.INJECT1_0 = "NO";
    defparam add_1706_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0110000) 
//

module \ArmPeripheral(axis_haddr=8'b0110000)  (Stepper_A_M0_c_0, \register_addr[0] , 
            debug_c_c, n34066, n3862, VCC_net, GND_net, Stepper_A_nFault_c, 
            \read_size[0] , n14114, n29712, n14493, n579, n14555, 
            prev_select, n32155, \read_size[2] , n30019, n34068, Stepper_A_M1_c_1, 
            n34069, \steps_reg[9] , \steps_reg[6] , \steps_reg[5] , 
            \steps_reg[3] , n34065, prev_step_clk, n34, step_clk, 
            n32142, n24, n32, n32_adj_1, prev_step_clk_adj_2, step_clk_adj_3, 
            n32144, limit_c_3, n22, n32_adj_4, prev_step_clk_adj_5, 
            step_clk_adj_6, n32145, n22_adj_7, n224, \register_addr[1] , 
            n32138, n34071, \databus[1] , Stepper_A_M2_c_2, n610, 
            \control_reg[3] , \databus[3] , n608, Stepper_A_Dir_c, \databus[5] , 
            Stepper_A_En_c, \databus[6] , \control_reg[7] , \databus[7] , 
            \div_factor_reg[5] , n32137, \div_factor_reg[6] , \div_factor_reg[9] , 
            \databus[9] , \databus[10] , \databus[11] , \databus[13] , 
            n32216, \databus[22] , \databus[23] , \databus[24] , \databus[25] , 
            \databus[26] , \databus[27] , \databus[28] , \databus[29] , 
            \databus[30] , \databus[31] , \databus[21] , \databus[20] , 
            \databus[19] , \databus[18] , \databus[17] , \databus[16] , 
            \databus[15] , \databus[14] , \databus[12] , \databus[8] , 
            \div_factor_reg[3] , int_step, read_value, n9496, n7376, 
            n21455, n21447, n29759, n8594, n29758, n28061) /* synthesis syn_module_defined=1 */ ;
    output Stepper_A_M0_c_0;
    input \register_addr[0] ;
    input debug_c_c;
    input n34066;
    input [31:0]n3862;
    input VCC_net;
    input GND_net;
    input Stepper_A_nFault_c;
    output \read_size[0] ;
    input n14114;
    input n29712;
    input n14493;
    input n579;
    input n14555;
    output prev_select;
    input n32155;
    output \read_size[2] ;
    input n30019;
    input n34068;
    output Stepper_A_M1_c_1;
    input n34069;
    output \steps_reg[9] ;
    output \steps_reg[6] ;
    output \steps_reg[5] ;
    output \steps_reg[3] ;
    input n34065;
    input prev_step_clk;
    input n34;
    input step_clk;
    output n32142;
    output n24;
    input n32;
    input n32_adj_1;
    input prev_step_clk_adj_2;
    input step_clk_adj_3;
    output n32144;
    input limit_c_3;
    output n22;
    input n32_adj_4;
    input prev_step_clk_adj_5;
    input step_clk_adj_6;
    output n32145;
    output n22_adj_7;
    output [31:0]n224;
    input \register_addr[1] ;
    input n32138;
    input n34071;
    input \databus[1] ;
    output Stepper_A_M2_c_2;
    input n610;
    output \control_reg[3] ;
    input \databus[3] ;
    input n608;
    output Stepper_A_Dir_c;
    input \databus[5] ;
    output Stepper_A_En_c;
    input \databus[6] ;
    output \control_reg[7] ;
    input \databus[7] ;
    output \div_factor_reg[5] ;
    input n32137;
    output \div_factor_reg[6] ;
    output \div_factor_reg[9] ;
    input \databus[9] ;
    input \databus[10] ;
    input \databus[11] ;
    input \databus[13] ;
    input n32216;
    input \databus[22] ;
    input \databus[23] ;
    input \databus[24] ;
    input \databus[25] ;
    input \databus[26] ;
    input \databus[27] ;
    input \databus[28] ;
    input \databus[29] ;
    input \databus[30] ;
    input \databus[31] ;
    input \databus[21] ;
    input \databus[20] ;
    input \databus[19] ;
    input \databus[18] ;
    input \databus[17] ;
    input \databus[16] ;
    input \databus[15] ;
    input \databus[14] ;
    input \databus[12] ;
    input \databus[8] ;
    output \div_factor_reg[3] ;
    output int_step;
    output [31:0]read_value;
    input n9496;
    input n7376;
    input n21455;
    input n21447;
    input n29759;
    input n8594;
    input n29758;
    output n28061;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire limit_latched, n30354;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n30355, fault_latched, prev_step_clk_c, step_clk_c, n182, 
        prev_limit_latched, n30360, n30361, n30411, n30412, n30413, 
        n11159, n32143, n22_c, n27478, n27477, n27476, n27475, 
        n27474, n27473, n27472, n27471, n27470, n27469, n27468, 
        n27467, n27466, n27465, n27464;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [7:0]n8593;
    
    wire n27463;
    wire [31:0]n7311;
    
    wire n30356, n30362;
    wire [31:0]n7347;
    
    wire n29766, n29767, n29761, n29764, n29760, n29769, n29768, 
        n29765, n29770, n29763, n29762, n29771, n29772, n29773, 
        n29774, n29775, n29776, n29777, n29778, n29779, n29780, 
        n29781, n29782, n49, n62, n58, n50, n41, n60, n54, 
        n42, n52, n38, n56, n46;
    
    LUT4 i22851_3_lut (.A(Stepper_A_M0_c_0), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n30354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22851_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i0 (.D(n3862[0]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    LUT4 i22852_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n30355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22852_3_lut.init = 16'hcaca;
    IFS1P3DX fault_latched_178 (.D(Stepper_A_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n29712), .SP(n14114), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n14493), .CK(debug_c_c), .Q(Stepper_A_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk_c), .CK(debug_c_c), .Q(prev_step_clk_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n14555), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n32155), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n30019), .SP(n14114), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3862[31]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    LUT4 i22857_3_lut (.A(Stepper_A_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n30360)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22857_3_lut.init = 16'hcaca;
    LUT4 i22858_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n30361)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22858_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i30 (.D(n3862[30]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3862[29]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3862[28]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3862[27]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3862[26]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3862[25]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3862[24]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3862[23]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3862[22]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3862[21]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3862[20]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3862[19]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3862[18]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3862[17]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3862[16]), .CK(debug_c_c), .CD(n34068), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3862[15]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3862[14]), .CK(debug_c_c), .CD(n34069), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3862[13]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3862[12]), .CK(debug_c_c), .CD(n34069), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3862[11]), .CK(debug_c_c), .CD(n34069), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3862[10]), .CK(debug_c_c), .CD(n34069), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3862[9]), .CK(debug_c_c), .CD(n34069), 
            .Q(\steps_reg[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3862[8]), .CK(debug_c_c), .CD(n34069), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3862[7]), .CK(debug_c_c), .CD(n34069), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3862[6]), .CK(debug_c_c), .CD(n34069), 
            .Q(\steps_reg[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3862[5]), .CK(debug_c_c), .CD(n34066), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3862[4]), .CK(debug_c_c), .CD(n34069), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3862[3]), .CK(debug_c_c), .CD(n34066), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3862[2]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3862[1]), .CK(debug_c_c), .CD(n34066), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    PFUMX i22910 (.BLUT(n30411), .ALUT(n30412), .C0(\register_addr[0] ), 
          .Z(n30413));
    LUT4 i4443_3_lut (.A(prev_limit_latched), .B(n34065), .C(limit_latched), 
         .Z(n11159)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i4443_3_lut.init = 16'hdcdc;
    LUT4 i2_3_lut_rep_321 (.A(prev_step_clk), .B(n34), .C(step_clk), .Z(n32142)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_321.init = 16'h4040;
    LUT4 i1_4_lut_4_lut (.A(prev_step_clk), .B(n34), .C(step_clk), .D(n34065), 
         .Z(n24)) /* synthesis lut_function=(!(A (C+(D))+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut.init = 16'h004a;
    LUT4 i2_3_lut_rep_322 (.A(n32), .B(prev_step_clk_c), .C(step_clk_c), 
         .Z(n32143)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_322.init = 16'h2020;
    LUT4 i1_4_lut_4_lut_adj_1 (.A(n32), .B(prev_step_clk_c), .C(step_clk_c), 
         .D(n34065), .Z(n22_c)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_1.init = 16'h002c;
    LUT4 i2_3_lut_rep_323 (.A(n32_adj_1), .B(prev_step_clk_adj_2), .C(step_clk_adj_3), 
         .Z(n32144)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_323.init = 16'h2020;
    LUT4 i118_1_lut (.A(limit_c_3), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_4_lut_adj_2 (.A(n32_adj_1), .B(prev_step_clk_adj_2), .C(step_clk_adj_3), 
         .D(n34065), .Z(n22)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_2.init = 16'h002c;
    LUT4 i2_3_lut_rep_324 (.A(n32_adj_4), .B(prev_step_clk_adj_5), .C(step_clk_adj_6), 
         .Z(n32145)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i2_3_lut_rep_324.init = 16'h2020;
    LUT4 i1_4_lut_4_lut_adj_3 (.A(n32_adj_4), .B(prev_step_clk_adj_5), .C(step_clk_adj_6), 
         .D(n34065), .Z(n22_adj_7)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(41[20:26])
    defparam i1_4_lut_4_lut_adj_3.init = 16'h002c;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27478), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27477), .COUT(n27478), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27476), .COUT(n27477), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27475), .COUT(n27476), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27474), .COUT(n27475), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27473), .COUT(n27474), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27472), .COUT(n27473), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27471), .COUT(n27472), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27470), .COUT(n27471), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27469), .COUT(n27470), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27468), .COUT(n27469), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(\steps_reg[9] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27467), .COUT(n27468), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27466), .COUT(n27467), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27465), .COUT(n27466), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27464), .COUT(n27465), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    LUT4 i15172_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n8593[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i15172_2_lut.init = 16'h2222;
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27463), .COUT(n27464), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    LUT4 mux_1990_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n7311[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1990_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1990_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n7311[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1990_i8_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(n32), .C1(step_clk_c), .D1(prev_step_clk_c), 
          .COUT(n27463), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    PFUMX i22853 (.BLUT(n30354), .ALUT(n30355), .C0(\register_addr[1] ), 
          .Z(n30356));
    PFUMX i22859 (.BLUT(n30360), .ALUT(n30361), .C0(\register_addr[1] ), 
          .Z(n30362));
    FD1P3JX control_reg_i2 (.D(\databus[1] ), .SP(n32138), .PD(n34071), 
            .CK(debug_c_c), .Q(Stepper_A_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n14493), .CK(debug_c_c), .Q(Stepper_A_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(\databus[3] ), .SP(n32138), .PD(n34071), 
            .CK(debug_c_c), .Q(\control_reg[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n14493), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(\databus[5] ), .SP(n32138), .PD(n34071), 
            .CK(debug_c_c), .Q(Stepper_A_Dir_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(\databus[6] ), .SP(n32138), .PD(n34071), 
            .CK(debug_c_c), .Q(Stepper_A_En_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(\databus[7] ), .SP(n32138), .CD(n11159), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n14555), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n14555), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(\databus[5] ), .SP(n32137), .PD(n34071), 
            .CK(debug_c_c), .Q(\div_factor_reg[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(\databus[6] ), .SP(n32137), .PD(n34071), 
            .CK(debug_c_c), .Q(\div_factor_reg[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(\databus[7] ), .SP(n32137), .PD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(\databus[9] ), .SP(n32137), .PD(n34071), 
            .CK(debug_c_c), .Q(\div_factor_reg[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(\databus[10] ), .SP(n32137), .PD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(\databus[11] ), .SP(n32137), .PD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(\databus[13] ), .SP(n32137), .PD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(\databus[22] ), .SP(n32137), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(\databus[23] ), .SP(n32137), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(\databus[24] ), .SP(n32137), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(\databus[25] ), .SP(n32137), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(\databus[26] ), .SP(n32137), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(\databus[27] ), .SP(n32137), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(\databus[28] ), .SP(n32137), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(\databus[29] ), .SP(n32137), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(\databus[30] ), .SP(n32137), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(\databus[31] ), .SP(n32137), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(\databus[21] ), .SP(n14555), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(\databus[20] ), .SP(n14555), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(\databus[19] ), .SP(n14555), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(\databus[18] ), .SP(n14555), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(\databus[17] ), .SP(n14555), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(\databus[16] ), .SP(n14555), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(\databus[15] ), .SP(n14555), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(\databus[14] ), .SP(n14555), .CD(n32216), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(\databus[12] ), .SP(n14555), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(\databus[8] ), .SP(n14555), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(\databus[3] ), .SP(n14555), .CD(n34071), 
            .CK(debug_c_c), .Q(\div_factor_reg[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(\databus[1] ), .SP(n14555), .CD(n34071), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3AX int_step_182 (.D(n32143), .SP(n22_c), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n30356), .SP(n14114), .CD(n9496), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30362), .SP(n14114), .CD(n9496), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30413), .SP(n14114), .CD(n9496), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n7376), .SP(n14114), .CD(n9496), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n7347[4]), .SP(n14114), .CD(n9496), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n21455), .SP(n14114), .CD(n9496), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n21447), .SP(n14114), .CD(n9496), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n7347[7]), .SP(n14114), .CD(n9496), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n29766), .SP(n14114), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n29759), .SP(n14114), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n29767), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n29761), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n29764), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n29760), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n29769), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n29768), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n29765), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n29770), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n29763), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n29762), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n29771), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n29772), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n29773), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n29774), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n29775), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n29776), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n29777), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n29778), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n29779), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n29780), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n29781), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n29782), .SP(n14114), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=625, LSE_RLINE=638 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    PFUMX mux_1994_i5 (.BLUT(n8593[4]), .ALUT(n7311[4]), .C0(\register_addr[1] ), 
          .Z(n7347[4]));
    PFUMX mux_1994_i8 (.BLUT(n8594), .ALUT(n7311[7]), .C0(\register_addr[1] ), 
          .Z(n7347[7]));
    LUT4 i1_4_lut (.A(div_factor_reg[8]), .B(n29758), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n29766)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_4 (.A(div_factor_reg[10]), .B(n29758), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n29767)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_4.init = 16'hc088;
    LUT4 i1_4_lut_adj_5 (.A(div_factor_reg[11]), .B(n29758), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n29761)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_5.init = 16'hc088;
    LUT4 i1_4_lut_adj_6 (.A(div_factor_reg[12]), .B(n29758), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n29764)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_6.init = 16'hc088;
    LUT4 i22908_3_lut (.A(Stepper_A_M2_c_2), .B(div_factor_reg[2]), .C(\register_addr[1] ), 
         .Z(n30411)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22908_3_lut.init = 16'hcaca;
    LUT4 i22909_3_lut (.A(n32), .B(steps_reg[2]), .C(\register_addr[1] ), 
         .Z(n30412)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22909_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_7 (.A(div_factor_reg[13]), .B(n29758), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n29760)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_7.init = 16'hc088;
    LUT4 i1_4_lut_adj_8 (.A(div_factor_reg[14]), .B(n29758), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n29769)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_8.init = 16'hc088;
    LUT4 i1_4_lut_adj_9 (.A(div_factor_reg[15]), .B(n29758), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n29768)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_9.init = 16'hc088;
    LUT4 i1_4_lut_adj_10 (.A(div_factor_reg[16]), .B(n29758), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n29765)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_10.init = 16'hc088;
    LUT4 i1_4_lut_adj_11 (.A(div_factor_reg[17]), .B(n29758), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n29770)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_11.init = 16'hc088;
    LUT4 i1_4_lut_adj_12 (.A(div_factor_reg[18]), .B(n29758), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n29763)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_12.init = 16'hc088;
    LUT4 i1_4_lut_adj_13 (.A(div_factor_reg[19]), .B(n29758), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n29762)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_13.init = 16'hc088;
    LUT4 i1_4_lut_adj_14 (.A(div_factor_reg[20]), .B(n29758), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n29771)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_14.init = 16'hc088;
    LUT4 i1_4_lut_adj_15 (.A(div_factor_reg[21]), .B(n29758), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n29772)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_15.init = 16'hc088;
    LUT4 i1_4_lut_adj_16 (.A(div_factor_reg[22]), .B(n29758), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n29773)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_16.init = 16'hc088;
    LUT4 i1_4_lut_adj_17 (.A(div_factor_reg[23]), .B(n29758), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n29774)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_17.init = 16'hc088;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n28061)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_18 (.A(div_factor_reg[24]), .B(n29758), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n29775)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_18.init = 16'hc088;
    LUT4 i1_4_lut_adj_19 (.A(div_factor_reg[25]), .B(n29758), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n29776)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_19.init = 16'hc088;
    LUT4 i1_4_lut_adj_20 (.A(div_factor_reg[26]), .B(n29758), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n29777)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_20.init = 16'hc088;
    LUT4 i1_4_lut_adj_21 (.A(div_factor_reg[27]), .B(n29758), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n29778)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_21.init = 16'hc088;
    LUT4 i1_4_lut_adj_22 (.A(div_factor_reg[28]), .B(n29758), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n29779)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_22.init = 16'hc088;
    LUT4 i17_4_lut (.A(steps_reg[21]), .B(steps_reg[27]), .C(steps_reg[15]), 
         .D(steps_reg[0]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[23]), .B(n52), .C(n38), .D(steps_reg[18]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[14]), .B(steps_reg[31]), .C(steps_reg[19]), 
         .D(steps_reg[11]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[7]), .B(\steps_reg[5] ), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[26]), .B(n56), .C(n46), .D(steps_reg[29]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[25]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_23 (.A(div_factor_reg[29]), .B(n29758), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n29780)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_23.init = 16'hc088;
    LUT4 i1_4_lut_adj_24 (.A(div_factor_reg[30]), .B(n29758), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n29781)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_24.init = 16'hc088;
    LUT4 i1_4_lut_adj_25 (.A(div_factor_reg[31]), .B(n29758), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n29782)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_25.init = 16'hc088;
    LUT4 i10_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[10]), .B(steps_reg[22]), .C(steps_reg[20]), 
         .D(\steps_reg[6] ), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(\steps_reg[9] ), .B(\steps_reg[3] ), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[28]), .C(steps_reg[13]), 
         .D(steps_reg[30]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[2]), .B(steps_reg[8]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    ClockDivider_U9 step_clk_gen (.n34065(n34065), .GND_net(GND_net), .div_factor_reg({div_factor_reg[31:10], 
            \div_factor_reg[9] , div_factor_reg[8:7], \div_factor_reg[6] , 
            \div_factor_reg[5] , div_factor_reg[4], \div_factor_reg[3] , 
            div_factor_reg[2:0]}), .step_clk(step_clk_c), .debug_c_c(debug_c_c), 
            .n34071(n34071)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U9
//

module ClockDivider_U9 (n34065, GND_net, div_factor_reg, step_clk, debug_c_c, 
            n34071) /* synthesis syn_module_defined=1 */ ;
    input n34065;
    input GND_net;
    input [31:0]div_factor_reg;
    output step_clk;
    input debug_c_c;
    input n34071;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[13:22])
    
    wire n8308, n32133;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n27151, n27150;
    wire [31:0]n40;
    
    wire n27390, n8342, n27389, n27149, n27148, n27388, n27387, 
        n27386, n27147, n27385, n27384, n27383, n27382, n27381, 
        n27380, n27379, n27146, n27378, n27145, n27377, n27144, 
        n27376, n27375, n8273, n16837, n27614;
    wire [31:0]n134;
    
    wire n27613, n27612, n27611, n27610, n27609, n27608, n27607, 
        n27606, n27143, n27605, n27604, n27603, n27602, n27601, 
        n27600, n27599, n27142, n27141, n27140, n27139, n27138, 
        n27137, n27136, n27135, n27166, n27165, n27164, n27163, 
        n27162, n27161, n27160, n27542, n27541, n27540, n27159, 
        n27539, n27538, n27537, n27536, n27535, n27534, n27533, 
        n27158, n27532, n27531, n27530, n27529, n27528, n27527, 
        n27157, n27156, n27155, n27154, n27153, n27152;
    
    LUT4 i1032_2_lut_rep_312 (.A(n8308), .B(n34065), .Z(n32133)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i1032_2_lut_rep_312.init = 16'heeee;
    CCU2D sub_2067_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27151));
    defparam sub_2067_add_2_1.INIT0 = 16'h0000;
    defparam sub_2067_add_2_1.INIT1 = 16'h5999;
    defparam sub_2067_add_2_1.INJECT1_0 = "NO";
    defparam sub_2067_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27150), .S1(n8308));
    defparam sub_2069_add_2_33.INIT0 = 16'h5999;
    defparam sub_2069_add_2_33.INIT1 = 16'h0000;
    defparam sub_2069_add_2_33.INJECT1_0 = "NO";
    defparam sub_2069_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27390), .S1(n8342));
    defparam sub_2070_add_2_33.INIT0 = 16'hf555;
    defparam sub_2070_add_2_33.INIT1 = 16'h0000;
    defparam sub_2070_add_2_33.INJECT1_0 = "NO";
    defparam sub_2070_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27389), .COUT(n27390));
    defparam sub_2070_add_2_31.INIT0 = 16'hf555;
    defparam sub_2070_add_2_31.INIT1 = 16'hf555;
    defparam sub_2070_add_2_31.INJECT1_0 = "NO";
    defparam sub_2070_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27149), .COUT(n27150));
    defparam sub_2069_add_2_31.INIT0 = 16'h5999;
    defparam sub_2069_add_2_31.INIT1 = 16'h5999;
    defparam sub_2069_add_2_31.INJECT1_0 = "NO";
    defparam sub_2069_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27148), .COUT(n27149));
    defparam sub_2069_add_2_29.INIT0 = 16'h5999;
    defparam sub_2069_add_2_29.INIT1 = 16'h5999;
    defparam sub_2069_add_2_29.INJECT1_0 = "NO";
    defparam sub_2069_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27388), .COUT(n27389));
    defparam sub_2070_add_2_29.INIT0 = 16'hf555;
    defparam sub_2070_add_2_29.INIT1 = 16'hf555;
    defparam sub_2070_add_2_29.INJECT1_0 = "NO";
    defparam sub_2070_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27387), .COUT(n27388));
    defparam sub_2070_add_2_27.INIT0 = 16'hf555;
    defparam sub_2070_add_2_27.INIT1 = 16'hf555;
    defparam sub_2070_add_2_27.INJECT1_0 = "NO";
    defparam sub_2070_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27386), .COUT(n27387));
    defparam sub_2070_add_2_25.INIT0 = 16'hf555;
    defparam sub_2070_add_2_25.INIT1 = 16'hf555;
    defparam sub_2070_add_2_25.INJECT1_0 = "NO";
    defparam sub_2070_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27147), .COUT(n27148));
    defparam sub_2069_add_2_27.INIT0 = 16'h5999;
    defparam sub_2069_add_2_27.INIT1 = 16'h5999;
    defparam sub_2069_add_2_27.INJECT1_0 = "NO";
    defparam sub_2069_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27385), .COUT(n27386));
    defparam sub_2070_add_2_23.INIT0 = 16'hf555;
    defparam sub_2070_add_2_23.INIT1 = 16'hf555;
    defparam sub_2070_add_2_23.INJECT1_0 = "NO";
    defparam sub_2070_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27384), .COUT(n27385));
    defparam sub_2070_add_2_21.INIT0 = 16'hf555;
    defparam sub_2070_add_2_21.INIT1 = 16'hf555;
    defparam sub_2070_add_2_21.INJECT1_0 = "NO";
    defparam sub_2070_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27383), .COUT(n27384));
    defparam sub_2070_add_2_19.INIT0 = 16'hf555;
    defparam sub_2070_add_2_19.INIT1 = 16'hf555;
    defparam sub_2070_add_2_19.INJECT1_0 = "NO";
    defparam sub_2070_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27382), .COUT(n27383));
    defparam sub_2070_add_2_17.INIT0 = 16'hf555;
    defparam sub_2070_add_2_17.INIT1 = 16'hf555;
    defparam sub_2070_add_2_17.INJECT1_0 = "NO";
    defparam sub_2070_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27381), .COUT(n27382));
    defparam sub_2070_add_2_15.INIT0 = 16'hf555;
    defparam sub_2070_add_2_15.INIT1 = 16'hf555;
    defparam sub_2070_add_2_15.INJECT1_0 = "NO";
    defparam sub_2070_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27380), .COUT(n27381));
    defparam sub_2070_add_2_13.INIT0 = 16'hf555;
    defparam sub_2070_add_2_13.INIT1 = 16'hf555;
    defparam sub_2070_add_2_13.INJECT1_0 = "NO";
    defparam sub_2070_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27379), .COUT(n27380));
    defparam sub_2070_add_2_11.INIT0 = 16'hf555;
    defparam sub_2070_add_2_11.INIT1 = 16'hf555;
    defparam sub_2070_add_2_11.INJECT1_0 = "NO";
    defparam sub_2070_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27146), .COUT(n27147));
    defparam sub_2069_add_2_25.INIT0 = 16'h5999;
    defparam sub_2069_add_2_25.INIT1 = 16'h5999;
    defparam sub_2069_add_2_25.INJECT1_0 = "NO";
    defparam sub_2069_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27378), .COUT(n27379));
    defparam sub_2070_add_2_9.INIT0 = 16'hf555;
    defparam sub_2070_add_2_9.INIT1 = 16'hf555;
    defparam sub_2070_add_2_9.INJECT1_0 = "NO";
    defparam sub_2070_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27145), .COUT(n27146));
    defparam sub_2069_add_2_23.INIT0 = 16'h5999;
    defparam sub_2069_add_2_23.INIT1 = 16'h5999;
    defparam sub_2069_add_2_23.INJECT1_0 = "NO";
    defparam sub_2069_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27377), .COUT(n27378));
    defparam sub_2070_add_2_7.INIT0 = 16'hf555;
    defparam sub_2070_add_2_7.INIT1 = 16'hf555;
    defparam sub_2070_add_2_7.INJECT1_0 = "NO";
    defparam sub_2070_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27144), .COUT(n27145));
    defparam sub_2069_add_2_21.INIT0 = 16'h5999;
    defparam sub_2069_add_2_21.INIT1 = 16'h5999;
    defparam sub_2069_add_2_21.INJECT1_0 = "NO";
    defparam sub_2069_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27376), .COUT(n27377));
    defparam sub_2070_add_2_5.INIT0 = 16'hf555;
    defparam sub_2070_add_2_5.INIT1 = 16'hf555;
    defparam sub_2070_add_2_5.INJECT1_0 = "NO";
    defparam sub_2070_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2070_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27375), .COUT(n27376));
    defparam sub_2070_add_2_3.INIT0 = 16'hf555;
    defparam sub_2070_add_2_3.INIT1 = 16'hf555;
    defparam sub_2070_add_2_3.INJECT1_0 = "NO";
    defparam sub_2070_add_2_3.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n8273), .CK(debug_c_c), .CD(n34071), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n32133), .PD(n16837), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    LUT4 i10145_2_lut_3_lut (.A(n8308), .B(n34065), .C(n8342), .Z(n16837)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i10145_2_lut_3_lut.init = 16'he0e0;
    CCU2D count_2665_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27614), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_33.INIT1 = 16'h0000;
    defparam count_2665_add_4_33.INJECT1_0 = "NO";
    defparam count_2665_add_4_33.INJECT1_1 = "NO";
    FD1S3IX count_2665__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i0.GSR = "ENABLED";
    CCU2D sub_2070_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27375));
    defparam sub_2070_add_2_1.INIT0 = 16'h0000;
    defparam sub_2070_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_2070_add_2_1.INJECT1_0 = "NO";
    defparam sub_2070_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27613), .COUT(n27614), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2665_add_4_31.INJECT1_0 = "NO";
    defparam count_2665_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27612), .COUT(n27613), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2665_add_4_29.INJECT1_0 = "NO";
    defparam count_2665_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27611), .COUT(n27612), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2665_add_4_27.INJECT1_0 = "NO";
    defparam count_2665_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27610), .COUT(n27611), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2665_add_4_25.INJECT1_0 = "NO";
    defparam count_2665_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27609), .COUT(n27610), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2665_add_4_23.INJECT1_0 = "NO";
    defparam count_2665_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27608), .COUT(n27609), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2665_add_4_21.INJECT1_0 = "NO";
    defparam count_2665_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27607), .COUT(n27608), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2665_add_4_19.INJECT1_0 = "NO";
    defparam count_2665_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27606), .COUT(n27607), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2665_add_4_17.INJECT1_0 = "NO";
    defparam count_2665_add_4_17.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27143), .COUT(n27144));
    defparam sub_2069_add_2_19.INIT0 = 16'h5999;
    defparam sub_2069_add_2_19.INIT1 = 16'h5999;
    defparam sub_2069_add_2_19.INJECT1_0 = "NO";
    defparam sub_2069_add_2_19.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27605), .COUT(n27606), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2665_add_4_15.INJECT1_0 = "NO";
    defparam count_2665_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27604), .COUT(n27605), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2665_add_4_13.INJECT1_0 = "NO";
    defparam count_2665_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27603), .COUT(n27604), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2665_add_4_11.INJECT1_0 = "NO";
    defparam count_2665_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27602), .COUT(n27603), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2665_add_4_9.INJECT1_0 = "NO";
    defparam count_2665_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27601), .COUT(n27602), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2665_add_4_7.INJECT1_0 = "NO";
    defparam count_2665_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27600), .COUT(n27601), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2665_add_4_5.INJECT1_0 = "NO";
    defparam count_2665_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27599), .COUT(n27600), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2665_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2665_add_4_3.INJECT1_0 = "NO";
    defparam count_2665_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2665_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27599), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665_add_4_1.INIT0 = 16'hF000;
    defparam count_2665_add_4_1.INIT1 = 16'h0555;
    defparam count_2665_add_4_1.INJECT1_0 = "NO";
    defparam count_2665_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27142), .COUT(n27143));
    defparam sub_2069_add_2_17.INIT0 = 16'h5999;
    defparam sub_2069_add_2_17.INIT1 = 16'h5999;
    defparam sub_2069_add_2_17.INJECT1_0 = "NO";
    defparam sub_2069_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27141), .COUT(n27142));
    defparam sub_2069_add_2_15.INIT0 = 16'h5999;
    defparam sub_2069_add_2_15.INIT1 = 16'h5999;
    defparam sub_2069_add_2_15.INJECT1_0 = "NO";
    defparam sub_2069_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27140), .COUT(n27141));
    defparam sub_2069_add_2_13.INIT0 = 16'h5999;
    defparam sub_2069_add_2_13.INIT1 = 16'h5999;
    defparam sub_2069_add_2_13.INJECT1_0 = "NO";
    defparam sub_2069_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27139), .COUT(n27140));
    defparam sub_2069_add_2_11.INIT0 = 16'h5999;
    defparam sub_2069_add_2_11.INIT1 = 16'h5999;
    defparam sub_2069_add_2_11.INJECT1_0 = "NO";
    defparam sub_2069_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27138), .COUT(n27139));
    defparam sub_2069_add_2_9.INIT0 = 16'h5999;
    defparam sub_2069_add_2_9.INIT1 = 16'h5999;
    defparam sub_2069_add_2_9.INJECT1_0 = "NO";
    defparam sub_2069_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27137), .COUT(n27138));
    defparam sub_2069_add_2_7.INIT0 = 16'h5999;
    defparam sub_2069_add_2_7.INIT1 = 16'h5999;
    defparam sub_2069_add_2_7.INJECT1_0 = "NO";
    defparam sub_2069_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27136), .COUT(n27137));
    defparam sub_2069_add_2_5.INIT0 = 16'h5999;
    defparam sub_2069_add_2_5.INIT1 = 16'h5999;
    defparam sub_2069_add_2_5.INJECT1_0 = "NO";
    defparam sub_2069_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27135), .COUT(n27136));
    defparam sub_2069_add_2_3.INIT0 = 16'h5999;
    defparam sub_2069_add_2_3.INIT1 = 16'h5999;
    defparam sub_2069_add_2_3.INJECT1_0 = "NO";
    defparam sub_2069_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_2069_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27135));
    defparam sub_2069_add_2_1.INIT0 = 16'h0000;
    defparam sub_2069_add_2_1.INIT1 = 16'h5999;
    defparam sub_2069_add_2_1.INJECT1_0 = "NO";
    defparam sub_2069_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n32133), .CD(n16837), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_2067_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27166), .S1(n8273));
    defparam sub_2067_add_2_33.INIT0 = 16'h5555;
    defparam sub_2067_add_2_33.INIT1 = 16'h0000;
    defparam sub_2067_add_2_33.INJECT1_0 = "NO";
    defparam sub_2067_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27165), .COUT(n27166));
    defparam sub_2067_add_2_31.INIT0 = 16'h5999;
    defparam sub_2067_add_2_31.INIT1 = 16'h5999;
    defparam sub_2067_add_2_31.INJECT1_0 = "NO";
    defparam sub_2067_add_2_31.INJECT1_1 = "NO";
    FD1S3IX count_2665__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i1.GSR = "ENABLED";
    CCU2D sub_2067_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27164), .COUT(n27165));
    defparam sub_2067_add_2_29.INIT0 = 16'h5999;
    defparam sub_2067_add_2_29.INIT1 = 16'h5999;
    defparam sub_2067_add_2_29.INJECT1_0 = "NO";
    defparam sub_2067_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27163), .COUT(n27164));
    defparam sub_2067_add_2_27.INIT0 = 16'h5999;
    defparam sub_2067_add_2_27.INIT1 = 16'h5999;
    defparam sub_2067_add_2_27.INJECT1_0 = "NO";
    defparam sub_2067_add_2_27.INJECT1_1 = "NO";
    FD1S3IX count_2665__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i2.GSR = "ENABLED";
    FD1S3IX count_2665__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i3.GSR = "ENABLED";
    FD1S3IX count_2665__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i4.GSR = "ENABLED";
    FD1S3IX count_2665__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i5.GSR = "ENABLED";
    FD1S3IX count_2665__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i6.GSR = "ENABLED";
    FD1S3IX count_2665__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i7.GSR = "ENABLED";
    FD1S3IX count_2665__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i8.GSR = "ENABLED";
    FD1S3IX count_2665__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i9.GSR = "ENABLED";
    FD1S3IX count_2665__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i10.GSR = "ENABLED";
    FD1S3IX count_2665__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i11.GSR = "ENABLED";
    FD1S3IX count_2665__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i12.GSR = "ENABLED";
    FD1S3IX count_2665__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i13.GSR = "ENABLED";
    FD1S3IX count_2665__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i14.GSR = "ENABLED";
    FD1S3IX count_2665__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i15.GSR = "ENABLED";
    FD1S3IX count_2665__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i16.GSR = "ENABLED";
    FD1S3IX count_2665__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i17.GSR = "ENABLED";
    FD1S3IX count_2665__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i18.GSR = "ENABLED";
    FD1S3IX count_2665__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i19.GSR = "ENABLED";
    FD1S3IX count_2665__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i20.GSR = "ENABLED";
    FD1S3IX count_2665__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i21.GSR = "ENABLED";
    FD1S3IX count_2665__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i22.GSR = "ENABLED";
    FD1S3IX count_2665__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i23.GSR = "ENABLED";
    FD1S3IX count_2665__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i24.GSR = "ENABLED";
    FD1S3IX count_2665__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i25.GSR = "ENABLED";
    FD1S3IX count_2665__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i26.GSR = "ENABLED";
    FD1S3IX count_2665__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i27.GSR = "ENABLED";
    FD1S3IX count_2665__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i28.GSR = "ENABLED";
    FD1S3IX count_2665__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i29.GSR = "ENABLED";
    FD1S3IX count_2665__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i30.GSR = "ENABLED";
    FD1S3IX count_2665__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n32133), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2665__i31.GSR = "ENABLED";
    CCU2D sub_2067_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27162), .COUT(n27163));
    defparam sub_2067_add_2_25.INIT0 = 16'h5999;
    defparam sub_2067_add_2_25.INIT1 = 16'h5999;
    defparam sub_2067_add_2_25.INJECT1_0 = "NO";
    defparam sub_2067_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27161), .COUT(n27162));
    defparam sub_2067_add_2_23.INIT0 = 16'h5999;
    defparam sub_2067_add_2_23.INIT1 = 16'h5999;
    defparam sub_2067_add_2_23.INJECT1_0 = "NO";
    defparam sub_2067_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27160), .COUT(n27161));
    defparam sub_2067_add_2_21.INIT0 = 16'h5999;
    defparam sub_2067_add_2_21.INIT1 = 16'h5999;
    defparam sub_2067_add_2_21.INJECT1_0 = "NO";
    defparam sub_2067_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27542), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27541), .COUT(n27542), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27540), .COUT(n27541), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27159), .COUT(n27160));
    defparam sub_2067_add_2_19.INIT0 = 16'h5999;
    defparam sub_2067_add_2_19.INIT1 = 16'h5999;
    defparam sub_2067_add_2_19.INJECT1_0 = "NO";
    defparam sub_2067_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27539), .COUT(n27540), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27538), .COUT(n27539), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27537), .COUT(n27538), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27536), .COUT(n27537), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27535), .COUT(n27536), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27534), .COUT(n27535), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27533), .COUT(n27534), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27158), .COUT(n27159));
    defparam sub_2067_add_2_17.INIT0 = 16'h5999;
    defparam sub_2067_add_2_17.INIT1 = 16'h5999;
    defparam sub_2067_add_2_17.INJECT1_0 = "NO";
    defparam sub_2067_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27532), .COUT(n27533), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27531), .COUT(n27532), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27530), .COUT(n27531), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27529), .COUT(n27530), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27528), .COUT(n27529), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27527), .COUT(n27528), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27527), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27157), .COUT(n27158));
    defparam sub_2067_add_2_15.INIT0 = 16'h5999;
    defparam sub_2067_add_2_15.INIT1 = 16'h5999;
    defparam sub_2067_add_2_15.INJECT1_0 = "NO";
    defparam sub_2067_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27156), .COUT(n27157));
    defparam sub_2067_add_2_13.INIT0 = 16'h5999;
    defparam sub_2067_add_2_13.INIT1 = 16'h5999;
    defparam sub_2067_add_2_13.INJECT1_0 = "NO";
    defparam sub_2067_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27155), .COUT(n27156));
    defparam sub_2067_add_2_11.INIT0 = 16'h5999;
    defparam sub_2067_add_2_11.INIT1 = 16'h5999;
    defparam sub_2067_add_2_11.INJECT1_0 = "NO";
    defparam sub_2067_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27154), .COUT(n27155));
    defparam sub_2067_add_2_9.INIT0 = 16'h5999;
    defparam sub_2067_add_2_9.INIT1 = 16'h5999;
    defparam sub_2067_add_2_9.INJECT1_0 = "NO";
    defparam sub_2067_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27153), .COUT(n27154));
    defparam sub_2067_add_2_7.INIT0 = 16'h5999;
    defparam sub_2067_add_2_7.INIT1 = 16'h5999;
    defparam sub_2067_add_2_7.INJECT1_0 = "NO";
    defparam sub_2067_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27152), .COUT(n27153));
    defparam sub_2067_add_2_5.INIT0 = 16'h5999;
    defparam sub_2067_add_2_5.INIT1 = 16'h5999;
    defparam sub_2067_add_2_5.INJECT1_0 = "NO";
    defparam sub_2067_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_2067_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27151), .COUT(n27152));
    defparam sub_2067_add_2_3.INIT0 = 16'h5999;
    defparam sub_2067_add_2_3.INIT1 = 16'h5999;
    defparam sub_2067_add_2_3.INJECT1_0 = "NO";
    defparam sub_2067_add_2_3.INJECT1_1 = "NO";
    
endmodule

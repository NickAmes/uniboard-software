// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.4.1.213
// Netlist written on Sat Jan 16 19:19:02 2016
//
// Verilog Description of module UniboardTop
//

module UniboardTop (uart_rx, uart_tx, status_led, clk_12MHz, Stepper_X_Step, 
            Stepper_X_Dir, Stepper_X_M0, Stepper_X_M1, Stepper_X_M2, 
            Stepper_X_En, Stepper_X_nFault, Stepper_Y_Step, Stepper_Y_Dir, 
            Stepper_Y_M0, Stepper_Y_M1, Stepper_Y_M2, Stepper_Y_En, 
            Stepper_Y_nFault, Stepper_Z_Step, Stepper_Z_Dir, Stepper_Z_M0, 
            Stepper_Z_M1, Stepper_Z_M2, Stepper_Z_En, Stepper_Z_nFault, 
            Stepper_A_Step, Stepper_A_Dir, Stepper_A_M0, Stepper_A_M1, 
            Stepper_A_M2, Stepper_A_En, Stepper_A_nFault, limit, expansion1, 
            expansion2, expansion3, expansion4, expansion5, signal_light, 
            encoder_ra, encoder_rb, encoder_ri, encoder_la, encoder_lb, 
            encoder_li, rc_ch1, rc_ch2, rc_ch3, rc_ch4, rc_ch7, 
            rc_ch8, motor_pwm_l, motor_pwm_r, xbee_pause, debug) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[8:19])
    input uart_rx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[13:20])
    output uart_tx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[14:21])
    output [2:0]status_led;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    input clk_12MHz;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    output Stepper_X_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:31])
    output Stepper_X_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:30])
    output Stepper_X_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    output Stepper_X_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    output Stepper_X_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    output Stepper_X_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[17:29])
    input Stepper_X_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(375[16:32])
    output Stepper_Y_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:31])
    output Stepper_Y_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:30])
    output Stepper_Y_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    output Stepper_Y_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    output Stepper_Y_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    output Stepper_Y_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[17:29])
    input Stepper_Y_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(383[16:32])
    output Stepper_Z_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:31])
    output Stepper_Z_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:30])
    output Stepper_Z_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    output Stepper_Z_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    output Stepper_Z_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    output Stepper_Z_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[17:29])
    input Stepper_Z_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(391[16:32])
    output Stepper_A_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:31])
    output Stepper_A_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:30])
    output Stepper_A_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    output Stepper_A_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    output Stepper_A_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    output Stepper_A_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[17:29])
    input Stepper_A_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(399[16:32])
    input [3:0]limit;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    output expansion1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    output expansion2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    output expansion3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[14:24])
    output expansion4 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    output expansion5 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[13:23])
    output signal_light;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(407[14:26])
    input encoder_ra;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    input encoder_rb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    input encoder_ri;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    input encoder_la;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    input encoder_lb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    input encoder_li;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(414[13:23])
    input rc_ch1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    input rc_ch2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    input rc_ch3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    input rc_ch4;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    input rc_ch7;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    input rc_ch8;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(421[13:19])
    output motor_pwm_l;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    output motor_pwm_r;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[14:25])
    input xbee_pause;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(425[13:23])
    output [8:0]debug;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [127:0]select /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    
    wire GND_net, VCC_net, n9388_c, n9387, Stepper_X_Step_c, Stepper_X_Dir_c, 
        Stepper_X_M0_c_0, Stepper_X_M1_c_1, Stepper_X_M2_c_2, Stepper_X_En_c, 
        Stepper_X_nFault_c, Stepper_Y_Step_c, Stepper_Y_Dir_c, Stepper_Y_M0_c_0, 
        Stepper_Y_M1_c_1, Stepper_Y_M2_c_2, Stepper_Y_En_c, Stepper_Y_nFault_c, 
        Stepper_Z_Step_c, Stepper_Z_Dir_c, Stepper_Z_M0_c_0, Stepper_Z_M1_c_1, 
        Stepper_Z_M2_c_2, Stepper_Z_En_c, Stepper_Z_nFault_c, Stepper_A_Step_c, 
        Stepper_A_Dir_c, Stepper_A_M0_c_0, Stepper_A_M1_c_1, Stepper_A_M2_c_2, 
        Stepper_A_En_c, Stepper_A_nFault_c, limit_c_3, limit_c_2, limit_c_1, 
        limit_c_0, signal_light_c, rc_ch1_c, rc_ch2_c, rc_ch3_c, rc_ch4_c, 
        rc_ch7_c, rc_ch8_c, xbee_pause_c, debug_c_7, debug_c_5, debug_c_4, 
        debug_c_3, debug_c_2;
    wire [31:0]databus;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(458[14:21])
    wire [2:0]reg_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(459[13:21])
    wire [7:0]register_addr;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    
    wire rw, n84, n24974, n12590;
    wire [15:0]reset_count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    
    wire n1, n13, n24988, n27575, n21, n28921;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    wire [31:0]databus_out;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(55[13:24])
    
    wire n27509, n27638, n2, n26342, n14286, n5, n18750, n28920;
    wire [31:0]n1286;
    
    wire n26939, n88, n1030, n27442, n12230, n19982, n27046, n28918, 
        n28917, n1_adj_389, n1_adj_390, n15;
    wire [31:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    wire [31:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(30[13:23])
    wire [2:0]read_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(31[12:21])
    
    wire n11908;
    wire [7:0]n7885;
    
    wire n60, n28914, n28913, n28912, n11618, n11636, n30, n4, 
        n28911, n14, n241;
    wire [7:0]read_value_adj_650;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(63[12:22])
    wire [2:0]read_size_adj_651;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(64[12:21])
    
    wire n64, n27556;
    wire [15:0]n281;
    
    wire n2_adj_399;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]read_value_adj_655;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_656;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select, n3359, n2_adj_434, n26778, n27050, n12104;
    wire [7:0]n572;
    
    wire n3446;
    wire [7:0]control_reg_adj_664;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]steps_reg_adj_666;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire stepping;
    wire [31:0]read_value_adj_667;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_668;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_470, n53, n1_adj_471, n6, n7904, n27079, 
        n10501, n28910, n24993;
    wire [7:0]n572_adj_684;
    
    wire n1_adj_472;
    wire [7:0]control_reg_adj_703;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]steps_reg_adj_705;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire stepping_adj_476;
    wire [31:0]read_value_adj_706;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_707;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_511, n27527, n3585, n3176, n12064, n6_adj_512, 
        n12042, motor_pwm_l_c;
    wire [7:0]control_reg_adj_742;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]div_factor_reg_adj_743;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg_adj_744;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire stepping_adj_516;
    wire [31:0]read_value_adj_745;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_746;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_551, n3582, n20503, n10489, n29063, n48, 
        n29056, n16, n12, n1_adj_552, n27033, n29052, n26917, 
        n11997, n11996, n10, n28905;
    wire [31:0]n581_adj_763;
    
    wire n1_adj_553, n28904, n176, n7844, n28903, n28901, n24991, 
        n24690, n14_adj_554, n27026, n30644, n27014, n15_adj_555, 
        n14_adj_556, n15_adj_557, n24994, n27444, n11947, n27443, 
        n14439, n26690, n27029, n4_adj_558, n15_adj_559, n28900, 
        n11, n10_adj_560, n9, n8, n28899, n30653, n2_adj_561, 
        n27025, n1_adj_562, n4_adj_563;
    wire [14:0]n66_adj_1089;
    
    wire n4_adj_564, n4_adj_565, n1_adj_566, n6_adj_567, n27640, n16_adj_568, 
        n14_adj_569, n12_adj_570, n10_adj_571, n8_adj_572, n6_adj_573, 
        n5_adj_574, n4_adj_575, n27040, n4_adj_576, n4_adj_577, n30652, 
        n1_adj_578, n2_adj_579, n1_adj_580, n2_adj_581, n1_adj_582, 
        n2_adj_583, n1_adj_584, n2_adj_585, n4_adj_586, n4_adj_587, 
        n1_adj_588, n2_adj_589, n1_adj_590, n2_adj_591, n1_adj_592, 
        n2_adj_593, n29028, n1_adj_594, n2_adj_595, n1_adj_596, n2_adj_597, 
        n1_adj_598, n2_adj_599, n1_adj_600, n2_adj_601, n29025, n1_adj_602, 
        n2_adj_603, n1_adj_604, n2_adj_605, n27582, n1_adj_606, n2_adj_607, 
        n29021, n24976, n7840, n2_adj_608, n8_adj_609, n6_adj_610, 
        n29018, n29016, n2_adj_611, n27080, n24911;
    wire [31:0]n6092;
    
    wire n27065, n29011, n27023, n29008, n6_adj_612, n14053, n28898, 
        n26918, n26915, n14_adj_613;
    wire [12:0]count_adj_802;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    wire [12:0]count_adj_805;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    wire [7:0]n7895;
    
    wire n26869, n28991, n28990, motor_pwm_r_c, n24442, n27024, 
        n27395, n2_adj_621, n24441, n26777, n4_adj_622, n28981, 
        n30651, n27081, n27387, n24440, n24439, n1_adj_623, n24438, 
        n27382, n28974, n28973, n24437, n28972, n12807, n7894, 
        n24436, n12804, n2_adj_624, n7, n28966, n8050, n8044, 
        n8040, n27493, n28965, n28964, n27372, n28960, n28959, 
        n28958, n14380, n28957, n14379, n28956, n28955, n27035, 
        n17, n30650, n27037, n26870, n27039, n27031, n27364, n27049, 
        n12754, n27045, n28888, n27048, n27034, n54, n25126, n27569, 
        n24998, n1_adj_625, n27028, n30649, n27030, n6670, n27359, 
        n28946, n27032, n27041, n27036, n1018, n27042, n27044, 
        n27043, n27038, n27027, n27047, n27590, n28937, n28936, 
        n28935, n27548, n28934, n28932, n2_adj_626, n30648, n2_adj_627, 
        n30647, n28931, n9_adj_628, n28893, n28929, n28928, n28927, 
        n24970, n22447, n11253;
    
    VHI i2 (.Z(VCC_net));
    PWMPeripheral motor_pwm (.\read_size[0] (read_size_adj_651[0]), .debug_c_c(debug_c_c), 
            .n28920(n28920), .n30649(n30649), .\databus[0] (databus[0]), 
            .\select[2] (select[2]), .n282(n281[15]), .n30653(n30653), 
            .\databus[6] (databus[6]), .\databus[5] (databus[5]), .\databus[4] (databus[4]), 
            .\databus[3] (databus[3]), .\databus[2] (databus[2]), .\databus[1] (databus[1]), 
            .n29063(n29063), .n28900(n28900), .n30647(n30647), .\register_addr[0] (register_addr[0]), 
            .rw(rw), .read_value({read_value_adj_650}), .n8044(n8044), 
            .n64(n64), .\count[0] (count_adj_805[0]), .n10489(n10489), 
            .n28893(n28893), .GND_net(GND_net), .n7885({n7885}), .n7894(n7894), 
            .\count[3] (count_adj_805[3]), .n14286(n14286), .\count[7] (count_adj_805[7]), 
            .\count[5] (count_adj_805[5]), .\count[1] (count_adj_805[1]), 
            .\count[6] (count_adj_805[6]), .\count[8] (count_adj_805[8]), 
            .\count[4] (count_adj_805[4]), .\count[2] (count_adj_805[2]), 
            .motor_pwm_r_c(motor_pwm_r_c), .n3585(n3585), .\count[0]_adj_185 (count_adj_802[0]), 
            .n10501(n10501), .n14439(n14439), .\count[12] (count_adj_802[12]), 
            .\count[11] (count_adj_802[11]), .\count[9] (count_adj_802[9]), 
            .\count[8]_adj_186 (count_adj_802[8]), .\count[6]_adj_187 (count_adj_802[6]), 
            .\count[5]_adj_188 (count_adj_802[5]), .\count[3]_adj_189 (count_adj_802[3]), 
            .\count[2]_adj_190 (count_adj_802[2]), .\count[1]_adj_191 (count_adj_802[1]), 
            .n28911(n28911), .n10(n10_adj_571), .n12(n12_adj_570), .\reset_count[5] (reset_count[5]), 
            .n27079(n27079), .\reset_count[6] (reset_count[6]), .\reset_count[4] (reset_count[4]), 
            .n27080(n27080), .\reset_count[8] (reset_count[8]), .\reset_count[7] (reset_count[7]), 
            .n7904(n7904), .n7898(n7895[5]), .n7897(n7895[6]), .n7900(n7895[3]), 
            .n7902(n7895[1]), .n7901(n7895[2]), .n7903(n7895[0]), .motor_pwm_l_c(motor_pwm_l_c), 
            .n25126(n25126), .n28958(n28958), .n6(n6_adj_573), .n8(n8_adj_572), 
            .n3582(n3582), .n6_adj_192(n6_adj_512)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(512[16] 522[40])
    LUT4 i21073_3_lut (.A(div_factor_reg_adj_743[0]), .B(steps_reg_adj_744[0]), 
         .C(register_addr[0]), .Z(n27443)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21073_3_lut.init = 16'hcaca;
    LUT4 i21198_4_lut (.A(n4_adj_575), .B(n12_adj_570), .C(n28911), .D(n27364), 
         .Z(n14_adj_569)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i21198_4_lut.init = 16'hcacc;
    LUT4 i1_2_lut_rep_240_3_lut_4_lut (.A(n29025), .B(n28964), .C(n30644), 
         .D(prev_select), .Z(n28898)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_240_3_lut_4_lut.init = 16'h0004;
    LUT4 LessThan_1430_i4_4_lut (.A(count_adj_802[0]), .B(count_adj_802[1]), 
         .C(n7895[1]), .D(n7895[0]), .Z(n4_adj_575)) /* synthesis lut_function=(A (B+!(C))+!A !(B (C (D))+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1430_i4_4_lut.init = 16'h8ecf;
    LUT4 i21339_4_lut_rep_413 (.A(n27080), .B(reset_count[14]), .C(n26342), 
         .D(n19982), .Z(n30647)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam i21339_4_lut_rep_413.init = 16'h373f;
    LUT4 Select_3612_i4_2_lut_3_lut_4_lut (.A(n29025), .B(n28964), .C(read_value_adj_655[5]), 
         .D(n30644), .Z(n4_adj_577)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3612_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i21359_4_lut (.A(n28912), .B(n28911), .C(n28931), .D(n27359), 
         .Z(n27372)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i21359_4_lut.init = 16'habaa;
    LUT4 i20989_4_lut (.A(n28932), .B(n28958), .C(n28957), .D(n5_adj_574), 
         .Z(n27359)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i20989_4_lut.init = 16'h5554;
    LUT4 LessThan_1430_i5_2_lut (.A(n7895[2]), .B(count_adj_802[2]), .Z(n5_adj_574)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1430_i5_2_lut.init = 16'h6666;
    LUT4 Select_3611_i4_2_lut_3_lut_4_lut (.A(n29025), .B(n28964), .C(read_value_adj_655[6]), 
         .D(n30644), .Z(n4_adj_586)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3611_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3610_i4_2_lut_3_lut_4_lut (.A(n29025), .B(n28964), .C(read_value_adj_655[7]), 
         .D(rw), .Z(n4_adj_587)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3610_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3617_i4_2_lut_3_lut_4_lut (.A(n29025), .B(n28964), .C(read_value_adj_655[0]), 
         .D(rw), .Z(n4_adj_563)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3617_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3615_i4_2_lut_3_lut_4_lut (.A(n29025), .B(n28964), .C(read_value_adj_655[2]), 
         .D(rw), .Z(n4_adj_564)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3615_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3614_i4_2_lut_3_lut_4_lut (.A(n29025), .B(n28964), .C(read_value_adj_655[3]), 
         .D(rw), .Z(n4_adj_565)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3614_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3613_i4_2_lut_3_lut_4_lut (.A(n29025), .B(n28964), .C(read_value_adj_655[4]), 
         .D(rw), .Z(n4_adj_576)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3613_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i4_3_lut_4_lut (.A(n29025), .B(n28964), .C(n8), .D(read_size_adj_656[0]), 
         .Z(n11)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;
    defparam i4_3_lut_4_lut.init = 16'hf4f0;
    PFUMX i13008 (.BLUT(n18750), .ALUT(n15_adj_559), .C0(register_addr[0]), 
          .Z(n6092[4]));
    LUT4 i21339_4_lut_rep_414 (.A(n27080), .B(reset_count[14]), .C(n26342), 
         .D(n19982), .Z(n30648)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam i21339_4_lut_rep_414.init = 16'h373f;
    LUT4 i21339_4_lut_rep_415 (.A(n27080), .B(reset_count[14]), .C(n26342), 
         .D(n19982), .Z(n30649)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam i21339_4_lut_rep_415.init = 16'h373f;
    LUT4 i21339_4_lut_rep_416 (.A(n27080), .B(reset_count[14]), .C(n26342), 
         .D(n19982), .Z(n30650)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam i21339_4_lut_rep_416.init = 16'h373f;
    LUT4 i21339_4_lut_rep_417 (.A(n27080), .B(reset_count[14]), .C(n26342), 
         .D(n19982), .Z(n30651)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam i21339_4_lut_rep_417.init = 16'h373f;
    LUT4 LessThan_1430_i13_2_lut_rep_273 (.A(n7895[6]), .B(count_adj_802[6]), 
         .Z(n28931)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1430_i13_2_lut_rep_273.init = 16'h6666;
    LUT4 LessThan_1430_i10_3_lut_3_lut (.A(n7895[6]), .B(count_adj_802[6]), 
         .C(count_adj_802[5]), .Z(n10_adj_571)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1430_i10_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i14099_2_lut_2_lut (.A(n30647), .B(databus[7]), .Z(n281[15])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14099_2_lut_2_lut.init = 16'h4444;
    LUT4 LessThan_1430_i11_2_lut_rep_274 (.A(n7895[5]), .B(count_adj_802[5]), 
         .Z(n28932)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1430_i11_2_lut_rep_274.init = 16'h6666;
    LUT4 i20994_2_lut_3_lut_4_lut (.A(n7895[5]), .B(count_adj_802[5]), .C(count_adj_802[6]), 
         .D(n7895[6]), .Z(n27364)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i20994_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i21339_4_lut_rep_418 (.A(n27080), .B(reset_count[14]), .C(n26342), 
         .D(n19982), .Z(n30652)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam i21339_4_lut_rep_418.init = 16'h373f;
    LUT4 i21339_4_lut_rep_419 (.A(n27080), .B(reset_count[14]), .C(n26342), 
         .D(n19982), .Z(n30653)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam i21339_4_lut_rep_419.init = 16'h373f;
    LUT4 LessThan_1433_i13_2_lut_rep_276 (.A(n7885[6]), .B(count_adj_805[6]), 
         .Z(n28934)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1433_i13_2_lut_rep_276.init = 16'h6666;
    LUT4 LessThan_1433_i10_3_lut_3_lut (.A(n7885[6]), .B(count_adj_805[6]), 
         .C(count_adj_805[5]), .Z(n10)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1433_i10_3_lut_3_lut.init = 16'hd4d4;
    LUT4 LessThan_1433_i11_2_lut_rep_277 (.A(n7885[5]), .B(count_adj_805[5]), 
         .Z(n28935)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1433_i11_2_lut_rep_277.init = 16'h6666;
    LUT4 i21017_2_lut_3_lut_4_lut (.A(n7885[5]), .B(count_adj_805[5]), .C(count_adj_805[6]), 
         .D(n7885[6]), .Z(n27387)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i21017_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 LessThan_1430_i17_2_lut_rep_254 (.A(n7904), .B(count_adj_802[8]), 
         .Z(n28912)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1430_i17_2_lut_rep_254.init = 16'h6666;
    LUT4 LessThan_1430_i16_3_lut_3_lut (.A(n7904), .B(count_adj_802[8]), 
         .C(n8_adj_572), .Z(n16_adj_568)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1430_i16_3_lut_3_lut.init = 16'hd4d4;
    LUT4 LessThan_1433_i15_2_lut_rep_255 (.A(n7885[7]), .B(count_adj_805[7]), 
         .Z(n28913)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1433_i15_2_lut_rep_255.init = 16'h6666;
    LUT4 i21230_4_lut (.A(n27081), .B(reset_count[14]), .C(n26342), .D(n19982), 
         .Z(n30)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam i21230_4_lut.init = 16'h373f;
    LUT4 i1_4_lut (.A(n20503), .B(n27079), .C(reset_count[6]), .D(reset_count[5]), 
         .Z(n27081)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[7:30])
    defparam i1_4_lut.init = 16'hfcec;
    LUT4 i14759_4_lut (.A(reset_count[0]), .B(reset_count[4]), .C(n6), 
         .D(reset_count[3]), .Z(n20503)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i14759_4_lut.init = 16'hccc8;
    LUT4 i2_2_lut (.A(reset_count[1]), .B(reset_count[2]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 LessThan_1433_i12_3_lut_3_lut (.A(n7885[7]), .B(count_adj_805[7]), 
         .C(n10), .Z(n12)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1433_i12_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i2_3_lut (.A(reset_count[12]), .B(reset_count[13]), .C(reset_count[11]), 
         .Z(n26342)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[7:30])
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i14252_2_lut (.A(reset_count[9]), .B(reset_count[10]), .Z(n19982)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14252_2_lut.init = 16'h8888;
    LUT4 LessThan_1433_i17_2_lut_rep_256 (.A(n7894), .B(count_adj_805[8]), 
         .Z(n28914)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1433_i17_2_lut_rep_256.init = 16'h6666;
    LUT4 i1_4_lut_adj_467 (.A(n19982), .B(reset_count[11]), .C(reset_count[8]), 
         .D(n24690), .Z(n26915)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_467.init = 16'h8880;
    FD1P3AX reset_count_2164_2165__i1 (.D(n66_adj_1089[0]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165__i1.GSR = "ENABLED";
    LUT4 LessThan_1433_i16_3_lut_3_lut (.A(n7894), .B(count_adj_805[8]), 
         .C(n8_adj_609), .Z(n16)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1433_i16_3_lut_3_lut.init = 16'hd4d4;
    LUT4 Select_3583_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[21]), 
         .D(n30644), .Z(n2_adj_607)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3583_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i21339_4_lut_rep_333 (.A(n27080), .B(reset_count[14]), .C(n26342), 
         .D(n19982), .Z(n28991)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam i21339_4_lut_rep_333.init = 16'h373f;
    LUT4 Select_3585_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[20]), 
         .D(rw), .Z(n2_adj_599)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3585_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3607_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[9]), 
         .D(rw), .Z(n2_adj_585)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3607_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n30647), .B(prev_select), .C(n28964), 
         .D(n29025), .Z(n11908)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h0010;
    PFUMX LessThan_1433_i18 (.BLUT(n14_adj_613), .ALUT(n16), .C0(n27395), 
          .Z(n3585));
    PFUMX i21074 (.BLUT(n27442), .ALUT(n27443), .C0(register_addr[1]), 
          .Z(n27444));
    LUT4 Select_3597_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[14]), 
         .D(n30644), .Z(n2_adj_593)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3597_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_241_3_lut_4_lut (.A(n28964), .B(n26939), .C(rw), 
         .D(prev_select_adj_511), .Z(n28899)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_241_3_lut_4_lut.init = 16'h0008;
    PFUMX LessThan_1430_i18 (.BLUT(n14_adj_569), .ALUT(n16_adj_568), .C0(n27372), 
          .Z(n3582));
    LUT4 i3_4_lut_rep_230 (.A(n54), .B(n6_adj_612), .C(n1030), .D(n4_adj_558), 
         .Z(n28888)) /* synthesis lut_function=(!(A ((C)+!B)+!A ((C+!(D))+!B))) */ ;
    defparam i3_4_lut_rep_230.init = 16'h0c08;
    LUT4 i13006_3_lut (.A(control_reg_adj_742[4]), .B(div_factor_reg_adj_743[4]), 
         .C(register_addr[1]), .Z(n18750)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13006_3_lut.init = 16'hcaca;
    LUT4 i21200_4_lut (.A(n4), .B(n12), .C(n28913), .D(n27387), .Z(n14_adj_613)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i21200_4_lut.init = 16'hcacc;
    LUT4 LessThan_1433_i4_4_lut (.A(count_adj_805[0]), .B(count_adj_805[1]), 
         .C(n7885[1]), .D(n7885[0]), .Z(n4)) /* synthesis lut_function=(A (B+!(C))+!A !(B (C (D))+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1433_i4_4_lut.init = 16'h8ecf;
    LUT4 i8385_2_lut_3_lut (.A(n54), .B(n6_adj_612), .C(n1030), .Z(n14053)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i8385_2_lut_3_lut.init = 16'h0808;
    IB xbee_pause_pad (.I(xbee_pause), .O(xbee_pause_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(425[13:23])
    IB rc_ch8_pad (.I(rc_ch8), .O(rc_ch8_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(421[13:19])
    IB rc_ch7_pad (.I(rc_ch7), .O(rc_ch7_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    IB rc_ch4_pad (.I(rc_ch4), .O(rc_ch4_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    IB rc_ch3_pad (.I(rc_ch3), .O(rc_ch3_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    IB rc_ch2_pad (.I(rc_ch2), .O(rc_ch2_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    IB rc_ch1_pad (.I(rc_ch1), .O(rc_ch1_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    IB limit_pad_0 (.I(limit[0]), .O(limit_c_0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_1 (.I(limit[1]), .O(limit_c_1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_2 (.I(limit[2]), .O(limit_c_2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_3 (.I(limit[3]), .O(limit_c_3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB Stepper_A_nFault_pad (.I(Stepper_A_nFault), .O(Stepper_A_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(399[16:32])
    IB Stepper_Z_nFault_pad (.I(Stepper_Z_nFault), .O(Stepper_Z_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(391[16:32])
    IB Stepper_Y_nFault_pad (.I(Stepper_Y_nFault), .O(Stepper_Y_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(383[16:32])
    IB Stepper_X_nFault_pad (.I(Stepper_X_nFault), .O(Stepper_X_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(375[16:32])
    IB debug_c_pad (.I(clk_12MHz), .O(debug_c_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    IB n9388_pad (.I(uart_rx), .O(n9388_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[13:20])
    OB debug_pad_0 (.I(n9388_c), .O(debug[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_1 (.I(n9387), .O(debug[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_2 (.I(debug_c_2), .O(debug[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_3 (.I(debug_c_3), .O(debug[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_4 (.I(debug_c_4), .O(debug[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_5 (.I(debug_c_5), .O(debug[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_6 (.I(n30647), .O(debug[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_7 (.I(debug_c_7), .O(debug[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_8 (.I(debug_c_c), .O(debug[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB motor_pwm_r_pad (.I(motor_pwm_r_c), .O(motor_pwm_r));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[14:25])
    OB motor_pwm_l_pad (.I(motor_pwm_l_c), .O(motor_pwm_l));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    OB signal_light_pad (.I(signal_light_c), .O(signal_light));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(407[14:26])
    OB expansion5_pad (.I(GND_net), .O(expansion5));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[13:23])
    OB expansion4_pad (.I(GND_net), .O(expansion4));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    OB expansion3_pad (.I(GND_net), .O(expansion3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[14:24])
    OB expansion2_pad (.I(GND_net), .O(expansion2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    OB expansion1_pad (.I(GND_net), .O(expansion1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    OB Stepper_A_En_pad (.I(Stepper_A_En_c), .O(Stepper_A_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[17:29])
    OB Stepper_A_M2_pad (.I(Stepper_A_M2_c_2), .O(Stepper_A_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    OB Stepper_A_M1_pad (.I(Stepper_A_M1_c_1), .O(Stepper_A_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    OB Stepper_A_M0_pad (.I(Stepper_A_M0_c_0), .O(Stepper_A_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    OB Stepper_A_Dir_pad (.I(Stepper_A_Dir_c), .O(Stepper_A_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:30])
    OB Stepper_A_Step_pad (.I(Stepper_A_Step_c), .O(Stepper_A_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:31])
    OB Stepper_Z_En_pad (.I(Stepper_Z_En_c), .O(Stepper_Z_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[17:29])
    OB Stepper_Z_M2_pad (.I(Stepper_Z_M2_c_2), .O(Stepper_Z_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    OB Stepper_Z_M1_pad (.I(Stepper_Z_M1_c_1), .O(Stepper_Z_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    OB Stepper_Z_M0_pad (.I(Stepper_Z_M0_c_0), .O(Stepper_Z_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    OB Stepper_Z_Dir_pad (.I(Stepper_Z_Dir_c), .O(Stepper_Z_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:30])
    OB Stepper_Z_Step_pad (.I(Stepper_Z_Step_c), .O(Stepper_Z_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:31])
    OB Stepper_Y_En_pad (.I(Stepper_Y_En_c), .O(Stepper_Y_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[17:29])
    OB Stepper_Y_M2_pad (.I(Stepper_Y_M2_c_2), .O(Stepper_Y_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    OB Stepper_Y_M1_pad (.I(Stepper_Y_M1_c_1), .O(Stepper_Y_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    OB Stepper_Y_M0_pad (.I(Stepper_Y_M0_c_0), .O(Stepper_Y_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    OB Stepper_Y_Dir_pad (.I(Stepper_Y_Dir_c), .O(Stepper_Y_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:30])
    OB Stepper_Y_Step_pad (.I(Stepper_Y_Step_c), .O(Stepper_Y_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:31])
    OB Stepper_X_En_pad (.I(Stepper_X_En_c), .O(Stepper_X_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[17:29])
    OB Stepper_X_M2_pad (.I(Stepper_X_M2_c_2), .O(Stepper_X_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    OB Stepper_X_M1_pad (.I(Stepper_X_M1_c_1), .O(Stepper_X_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    OB Stepper_X_M0_pad (.I(Stepper_X_M0_c_0), .O(Stepper_X_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    OB Stepper_X_Dir_pad (.I(Stepper_X_Dir_c), .O(Stepper_X_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:30])
    OB Stepper_X_Step_pad (.I(Stepper_X_Step_c), .O(Stepper_X_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:31])
    OB status_led_pad_0 (.I(VCC_net), .O(status_led[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    OB status_led_pad_1 (.I(VCC_net), .O(status_led[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    LUT4 i21351_4_lut (.A(n28914), .B(n28913), .C(n28934), .D(n27382), 
         .Z(n27395)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i21351_4_lut.init = 16'habaa;
    LUT4 i21012_4_lut (.A(n28935), .B(n28959), .C(n28960), .D(n5), .Z(n27382)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i21012_4_lut.init = 16'h5554;
    LUT4 LessThan_1433_i5_2_lut (.A(n7885[2]), .B(count_adj_805[2]), .Z(n5)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1433_i5_2_lut.init = 16'h6666;
    OB status_led_pad_2 (.I(VCC_net), .O(status_led[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    OB uart_tx_pad (.I(n9387), .O(uart_tx));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[14:21])
    LUT4 i21072_3_lut (.A(Stepper_A_M0_c_0), .B(stepping_adj_516), .C(register_addr[0]), 
         .Z(n27442)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21072_3_lut.init = 16'hcaca;
    LUT4 Select_3609_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[8]), 
         .D(n30644), .Z(n2_adj_581)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3609_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i14102_2_lut_2_lut (.A(n30647), .B(databus[6]), .Z(n572[6])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14102_2_lut_2_lut.init = 16'h4444;
    LUT4 i14200_2_lut_2_lut (.A(n30647), .B(databus[2]), .Z(n581_adj_763[2])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14200_2_lut_2_lut.init = 16'h4444;
    LUT4 i14205_2_lut_2_lut (.A(n30647), .B(databus[4]), .Z(n581_adj_763[4])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14205_2_lut_2_lut.init = 16'h4444;
    LUT4 i21260_4_lut_4_lut (.A(n28981), .B(n4_adj_622), .C(n9_adj_628), 
         .D(n1286[14]), .Z(n12064)) /* synthesis lut_function=(!((B (C+!(D))+!B !(D))+!A)) */ ;
    defparam i21260_4_lut_4_lut.init = 16'h2a00;
    FD1P3AX reset_count_2164_2165__i2 (.D(n66_adj_1089[1]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165__i2.GSR = "ENABLED";
    LUT4 i3_4_lut_4_lut (.A(n28981), .B(n1286[8]), .C(n29016), .D(n1286[0]), 
         .Z(n12754)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i3_4_lut_4_lut.init = 16'hfffd;
    LUT4 Select_3603_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[11]), 
         .D(n30644), .Z(n2_adj_583)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3603_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    CCU2D reset_count_2164_2165_add_4_15 (.A0(reset_count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n24442), .S0(n66_adj_1089[13]), 
          .S1(n66_adj_1089[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165_add_4_15.INIT0 = 16'hfaaa;
    defparam reset_count_2164_2165_add_4_15.INIT1 = 16'hfaaa;
    defparam reset_count_2164_2165_add_4_15.INJECT1_0 = "NO";
    defparam reset_count_2164_2165_add_4_15.INJECT1_1 = "NO";
    CCU2D reset_count_2164_2165_add_4_13 (.A0(reset_count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n24441), .COUT(n24442), .S0(n66_adj_1089[11]), 
          .S1(n66_adj_1089[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165_add_4_13.INIT0 = 16'hfaaa;
    defparam reset_count_2164_2165_add_4_13.INIT1 = 16'hfaaa;
    defparam reset_count_2164_2165_add_4_13.INJECT1_0 = "NO";
    defparam reset_count_2164_2165_add_4_13.INJECT1_1 = "NO";
    LUT4 Select_3605_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[10]), 
         .D(n30644), .Z(n2_adj_579)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3605_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    CCU2D reset_count_2164_2165_add_4_11 (.A0(reset_count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n24440), .COUT(n24441), .S0(n66_adj_1089[9]), 
          .S1(n66_adj_1089[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165_add_4_11.INIT0 = 16'hfaaa;
    defparam reset_count_2164_2165_add_4_11.INIT1 = 16'hfaaa;
    defparam reset_count_2164_2165_add_4_11.INJECT1_0 = "NO";
    defparam reset_count_2164_2165_add_4_11.INJECT1_1 = "NO";
    CCU2D reset_count_2164_2165_add_4_9 (.A0(reset_count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n24439), .COUT(n24440), .S0(n66_adj_1089[7]), 
          .S1(n66_adj_1089[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165_add_4_9.INIT0 = 16'hfaaa;
    defparam reset_count_2164_2165_add_4_9.INIT1 = 16'hfaaa;
    defparam reset_count_2164_2165_add_4_9.INJECT1_0 = "NO";
    defparam reset_count_2164_2165_add_4_9.INJECT1_1 = "NO";
    CCU2D reset_count_2164_2165_add_4_7 (.A0(reset_count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n24438), .COUT(n24439), .S0(n66_adj_1089[5]), 
          .S1(n66_adj_1089[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165_add_4_7.INIT0 = 16'hfaaa;
    defparam reset_count_2164_2165_add_4_7.INIT1 = 16'hfaaa;
    defparam reset_count_2164_2165_add_4_7.INJECT1_0 = "NO";
    defparam reset_count_2164_2165_add_4_7.INJECT1_1 = "NO";
    LUT4 Select_3601_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[12]), 
         .D(n30644), .Z(n2_adj_589)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3601_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3599_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[13]), 
         .D(n30644), .Z(n2_adj_591)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3599_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    CCU2D reset_count_2164_2165_add_4_5 (.A0(reset_count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n24437), .COUT(n24438), .S0(n66_adj_1089[3]), 
          .S1(n66_adj_1089[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165_add_4_5.INIT0 = 16'hfaaa;
    defparam reset_count_2164_2165_add_4_5.INIT1 = 16'hfaaa;
    defparam reset_count_2164_2165_add_4_5.INJECT1_0 = "NO";
    defparam reset_count_2164_2165_add_4_5.INJECT1_1 = "NO";
    CCU2D reset_count_2164_2165_add_4_3 (.A0(reset_count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n24436), .COUT(n24437), .S0(n66_adj_1089[1]), 
          .S1(n66_adj_1089[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165_add_4_3.INIT0 = 16'hfaaa;
    defparam reset_count_2164_2165_add_4_3.INIT1 = 16'hfaaa;
    defparam reset_count_2164_2165_add_4_3.INJECT1_0 = "NO";
    defparam reset_count_2164_2165_add_4_3.INJECT1_1 = "NO";
    CCU2D reset_count_2164_2165_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(reset_count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n24436), .S1(n66_adj_1089[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165_add_4_1.INIT0 = 16'hF000;
    defparam reset_count_2164_2165_add_4_1.INIT1 = 16'h0555;
    defparam reset_count_2164_2165_add_4_1.INJECT1_0 = "NO";
    defparam reset_count_2164_2165_add_4_1.INJECT1_1 = "NO";
    LUT4 Select_3595_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[15]), 
         .D(rw), .Z(n2_adj_603)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3595_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3593_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[16]), 
         .D(rw), .Z(n2_adj_605)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3593_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    GSR GSR_INST (.GSR(VCC_net));
    FD1P3AX reset_count_2164_2165__i3 (.D(n66_adj_1089[2]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165__i3.GSR = "ENABLED";
    FD1P3AX reset_count_2164_2165__i4 (.D(n66_adj_1089[3]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165__i4.GSR = "ENABLED";
    FD1P3AX reset_count_2164_2165__i5 (.D(n66_adj_1089[4]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165__i5.GSR = "ENABLED";
    FD1P3AX reset_count_2164_2165__i6 (.D(n66_adj_1089[5]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165__i6.GSR = "ENABLED";
    FD1P3AX reset_count_2164_2165__i7 (.D(n66_adj_1089[6]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165__i7.GSR = "ENABLED";
    FD1P3AX reset_count_2164_2165__i8 (.D(n66_adj_1089[7]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165__i8.GSR = "ENABLED";
    FD1P3AX reset_count_2164_2165__i9 (.D(n66_adj_1089[8]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165__i9.GSR = "ENABLED";
    FD1P3AX reset_count_2164_2165__i10 (.D(n66_adj_1089[9]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165__i10.GSR = "ENABLED";
    FD1P3AX reset_count_2164_2165__i11 (.D(n66_adj_1089[10]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165__i11.GSR = "ENABLED";
    FD1P3AX reset_count_2164_2165__i12 (.D(n66_adj_1089[11]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165__i12.GSR = "ENABLED";
    FD1P3AX reset_count_2164_2165__i13 (.D(n66_adj_1089[12]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165__i13.GSR = "ENABLED";
    FD1P3AX reset_count_2164_2165__i14 (.D(n66_adj_1089[13]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165__i14.GSR = "ENABLED";
    FD1P3AX reset_count_2164_2165__i15 (.D(n66_adj_1089[14]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2164_2165__i15.GSR = "ENABLED";
    LUT4 Select_3591_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[17]), 
         .D(rw), .Z(n2_adj_597)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3591_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3589_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[18]), 
         .D(rw), .Z(n2_adj_601)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3589_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3587_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[19]), 
         .D(rw), .Z(n2_adj_595)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3587_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    \ArmPeripheral(axis_haddr=8'b010000)  arm_y (.GND_net(GND_net), .n24974(n24974), 
            .stepping(stepping), .n14(n14_adj_556), .\register_addr[0] (register_addr[0]), 
            .n15(n15_adj_555), .\register_addr[1] (register_addr[1]), .Stepper_Y_M0_c_0(Stepper_Y_M0_c_0), 
            .debug_c_c(debug_c_c), .n30649(n30649), .VCC_net(VCC_net), 
            .Stepper_Y_nFault_c(Stepper_Y_nFault_c), .\read_size[0] (read_size_adj_668[0]), 
            .n26778(n26778), .n580(n572_adj_684[0]), .prev_select(prev_select_adj_470), 
            .n28974(n28974), .databus({databus}), .n3359(n3359), .n7840(n7840), 
            .n30651(n30651), .n30648(n30648), .n30650(n30650), .\control_reg[7] (control_reg_adj_664[7]), 
            .Stepper_Y_Dir_c(Stepper_Y_Dir_c), .n30652(n30652), .Stepper_Y_M2_c_2(Stepper_Y_M2_c_2), 
            .Stepper_Y_M1_c_1(Stepper_Y_M1_c_1), .\read_size[2] (read_size_adj_668[2]), 
            .n26869(n26869), .n30653(n30653), .\steps_reg[5] (steps_reg_adj_666[5]), 
            .\steps_reg[3] (steps_reg_adj_666[3]), .n30647(n30647), .Stepper_Y_En_c(Stepper_Y_En_c), 
            .Stepper_Y_Step_c(Stepper_Y_Step_c), .n8050(n8050), .read_value({read_value_adj_667}), 
            .n28966(n28966), .n28936(n28936), .\register_addr[5] (register_addr[5]), 
            .limit_c_1(limit_c_1), .n28991(n28991)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(574[25] 587[45])
    LUT4 LessThan_1430_i7_2_lut_rep_299 (.A(n7895[3]), .B(count_adj_802[3]), 
         .Z(n28957)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1430_i7_2_lut_rep_299.init = 16'h6666;
    \ProtocolInterface(baud_div=12)  protocol_interface (.n28973(n28973), 
            .n29056(n29056), .\read_value[22] (read_value_adj_745[22]), 
            .rw(rw), .n1(n1), .debug_c_c(debug_c_c), .n30644(n30644), 
            .n1318(n1286[0]), .register_addr({Open_0, Open_1, register_addr[5:4], 
            Open_2, Open_3, Open_4, Open_5}), .n29025(n29025), .debug_c_7(debug_c_7), 
            .\register_addr[1] (register_addr[1]), .\steps_reg[3] (steps_reg_adj_744[3]), 
            .n15(n15), .\register_addr[2] (register_addr[2]), .n28899(n28899), 
            .n28972(n28972), .n29008(n29008), .n7844(n7844), .n1304(n1286[14]), 
            .n1310(n1286[8]), .\register_addr[0] (register_addr[0]), .n12064(n12064), 
            .databus_out({databus_out}), .\read_value[21] (read_value_adj_745[21]), 
            .n1_adj_149(n1_adj_606), .n28921(n28921), .n12042(n12042), 
            .n8040(n8040), .databus({databus}), .\read_value[20] (read_value_adj_745[20]), 
            .n1_adj_150(n1_adj_598), .n9(n9_adj_628), .\sendcount[1] (sendcount[1]), 
            .\steps_reg[5] (steps_reg_adj_744[5]), .n14(n14), .n29052(n29052), 
            .n30647(n30647), .n12230(n12230), .\steps_reg[7] (steps_reg[7]), 
            .n13(n13), .n11636(n11636), .n28928(n28928), .n29011(n29011), 
            .n28990(n28990), .n11618(n11618), .prev_select(prev_select_adj_470), 
            .n28966(n28966), .n53(n53), .debug_c_2(debug_c_2), .\steps_reg[5]_adj_151 (steps_reg_adj_705[5]), 
            .n14_adj_152(n14_adj_554), .debug_c_3(debug_c_3), .debug_c_4(debug_c_4), 
            .debug_c_5(debug_c_5), .n28946(n28946), .prev_select_adj_153(prev_select_adj_551), 
            .n28910(n28910), .\read_value[16] (read_value_adj_745[16]), 
            .n1_adj_154(n1_adj_604), .\read_value[19] (read_value_adj_745[19]), 
            .n1_adj_155(n1_adj_594), .\read_value[15] (read_value_adj_745[15]), 
            .n1_adj_156(n1_adj_602), .\read_value[12] (read_value_adj_745[12]), 
            .n1_adj_157(n1_adj_588), .\read_value[13] (read_value_adj_745[13]), 
            .n1_adj_158(n1_adj_590), .\read_value[1] (read_value_adj_745[1]), 
            .n1_adj_159(n1_adj_566), .\read_value[18] (read_value_adj_745[18]), 
            .n1_adj_160(n1_adj_600), .\read_value[14] (read_value_adj_745[14]), 
            .n1_adj_161(n1_adj_592), .\read_value[17] (read_value_adj_745[17]), 
            .n1_adj_162(n1_adj_596), .n3359(n3359), .n28981(n28981), .\read_value[11] (read_value_adj_745[11]), 
            .n1_adj_163(n1_adj_582), .\read_value[10] (read_value_adj_745[10]), 
            .n1_adj_164(n1_adj_578), .\read_value[9] (read_value_adj_745[9]), 
            .n1_adj_165(n1_adj_584), .\read_value[8] (read_value_adj_745[8]), 
            .n1_adj_166(n1_adj_580), .\read_value[31] (read_value_adj_745[31]), 
            .n1_adj_167(n1_adj_562), .\read_value[30] (read_value_adj_745[30]), 
            .n1_adj_168(n1_adj_472), .\read_value[29] (read_value_adj_745[29]), 
            .n1_adj_169(n1_adj_552), .\read_value[28] (read_value_adj_745[28]), 
            .n1_adj_170(n1_adj_471), .\read_value[27] (read_value_adj_745[27]), 
            .n1_adj_171(n1_adj_389), .n22447(n22447), .\read_value[26] (read_value_adj_745[26]), 
            .n1_adj_172(n1_adj_390), .\read_value[25] (read_value_adj_745[25]), 
            .n1_adj_173(n1_adj_553), .\read_value[24] (read_value_adj_745[24]), 
            .n1_adj_174(n1_adj_623), .\steps_reg[3]_adj_175 (steps_reg_adj_705[3]), 
            .n15_adj_176(n15_adj_557), .\read_value[23] (read_value_adj_745[23]), 
            .n1_adj_177(n1_adj_625), .n26939(n26939), .n12590(n12590), 
            .n28929(n28929), .\select[4] (select[4]), .n28927(n28927), 
            .n29021(n29021), .n27014(n27014), .n14379(n14379), .n28937(n28937), 
            .n14380(n14380), .n3176(n3176), .n28974(n28974), .n26870(n26870), 
            .n26869(n26869), .n28917(n28917), .n28900(n28900), .n88(n88), 
            .n26777(n26777), .n26778(n26778), .n28964(n28964), .n28956(n28956), 
            .n28965(n28965), .\steps_reg[4] (steps_reg_adj_744[4]), .n15_adj_178(n15_adj_559), 
            .n29016(n29016), .n7840(n7840), .n48(n48), .\steps_reg[5]_adj_179 (steps_reg_adj_666[5]), 
            .n14_adj_180(n14_adj_556), .n84(n84), .\steps_reg[3]_adj_181 (steps_reg_adj_666[3]), 
            .n15_adj_182(n15_adj_555), .n60(n60), .n11253(n11253), .n11(n11), 
            .n9_adj_183(n9), .n10(n10_adj_560), .\reg_size[2] (reg_size[2]), 
            .n29018(n29018), .\select[1] (select[1]), .n12754(n12754), 
            .\select[2] (select[2]), .\select[7] (select[7]), .n28898(n28898), 
            .n3446(n3446), .n4(n4_adj_622), .n28936(n28936), .\reset_count[14] (reset_count[14]), 
            .n26915(n26915), .\reset_count[13] (reset_count[13]), .\reset_count[12] (reset_count[12]), 
            .\reset_count[7] (reset_count[7]), .\reset_count[6] (reset_count[6]), 
            .\reset_count[5] (reset_count[5]), .n24690(n24690), .n9387(n9387), 
            .GND_net(GND_net), .n9388_c(n9388_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(475[26] 485[57])
    LUT4 LessThan_1430_i6_3_lut_3_lut (.A(n7895[3]), .B(count_adj_802[3]), 
         .C(count_adj_802[2]), .Z(n6_adj_573)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1430_i6_3_lut_3_lut.init = 16'hd4d4;
    LUT4 LessThan_1433_i9_2_lut_rep_301 (.A(n7885[4]), .B(count_adj_805[4]), 
         .Z(n28959)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1433_i9_2_lut_rep_301.init = 16'h6666;
    LUT4 LessThan_1433_i8_3_lut_3_lut (.A(n7885[4]), .B(count_adj_805[4]), 
         .C(n6_adj_610), .Z(n8_adj_609)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1433_i8_3_lut_3_lut.init = 16'hd4d4;
    LUT4 LessThan_1433_i7_2_lut_rep_302 (.A(n7885[3]), .B(count_adj_805[3]), 
         .Z(n28960)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1433_i7_2_lut_rep_302.init = 16'h6666;
    LUT4 Select_3563_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[31]), 
         .D(n30644), .Z(n2_adj_561)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3563_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 LessThan_1433_i6_3_lut_3_lut (.A(n7885[3]), .B(count_adj_805[3]), 
         .C(count_adj_805[2]), .Z(n6_adj_610)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1433_i6_3_lut_3_lut.init = 16'hd4d4;
    LUT4 Select_3565_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[30]), 
         .D(rw), .Z(n2_adj_627)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3565_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i21_2_lut_rep_246_3_lut_4_lut (.A(select[4]), .B(n28990), .C(rw), 
         .D(n29025), .Z(n28904)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i21_2_lut_rep_246_3_lut_4_lut.init = 16'h0020;
    LUT4 Select_3567_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[29]), 
         .D(n30644), .Z(n2_adj_608)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3567_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    GlobalControlPeripheral global_control (.\select[1] (select[1]), .n30644(n30644), 
            .n29028(n29028), .rw(rw), .n6(n6_adj_567), .\read_value[2] (read_value[2]), 
            .debug_c_c(debug_c_c), .n12042(n12042), .n8040(n8040), .read_size({read_size}), 
            .n88(n88), .n30649(n30649), .signal_light_c(signal_light_c), 
            .n10501(n10501), .n14439(n14439), .\control_reg[7] (control_reg_adj_742[7]), 
            .n24911(n24911), .stepping(stepping_adj_516), .\control_reg[7]_adj_144 (control_reg[7]), 
            .n24994(n24994), .n21(n21), .\control_reg[7]_adj_145 (control_reg_adj_703[7]), 
            .n24970(n24970), .stepping_adj_146(stepping_adj_476), .n10489(n10489), 
            .n14286(n14286), .\control_reg[7]_adj_147 (control_reg_adj_664[7]), 
            .n24974(n24974), .stepping_adj_148(stepping), .\register[2][31] (\register[2] [31]), 
            .n30648(n30648), .\register[2][30] (\register[2] [30]), .\register[2][29] (\register[2] [29]), 
            .\register[2][28] (\register[2] [28]), .\register[2][27] (\register[2] [27]), 
            .\register[2][26] (\register[2] [26]), .\register[2][25] (\register[2] [25]), 
            .\register[2][24] (\register[2] [24]), .\register[2][23] (\register[2] [23]), 
            .\register[2][22] (\register[2] [22]), .\register[2][21] (\register[2] [21]), 
            .\register[2][20] (\register[2] [20]), .\register[2][19] (\register[2] [19]), 
            .\register[2][18] (\register[2] [18]), .\register[2][17] (\register[2] [17]), 
            .\register[2][16] (\register[2] [16]), .\register[2][15] (\register[2] [15]), 
            .\register[2][14] (\register[2] [14]), .\register[2][13] (\register[2] [13]), 
            .\register[2][12] (\register[2] [12]), .\register[2][11] (\register[2] [11]), 
            .\register[2][10] (\register[2] [10]), .\register[2][9] (\register[2] [9]), 
            .\register[2][8] (\register[2] [8]), .\register[2][7] (\register[2] [7]), 
            .\register[2][6] (\register[2] [6]), .\register[2][5] (\register[2] [5]), 
            .\register[2][4] (\register[2] [4]), .\register_addr[0] (register_addr[0]), 
            .n30647(n30647), .n28991(n28991), .xbee_pause_c(xbee_pause_c), 
            .\register_addr[5] (register_addr[5]), .n28972(n28972), .\register_addr[1] (register_addr[1]), 
            .\register_addr[2] (register_addr[2]), .n28920(n28920), .n22447(n22447), 
            .GND_net(GND_net), .n28921(n28921), .n29063(n29063), .n8044(n8044), 
            .n29025(n29025), .n29011(n29011), .n28901(n28901), .\read_value[3] (read_value[3]), 
            .\read_value[4] (read_value[4]), .n27030(n27030), .\read_value[5] (read_value[5]), 
            .n27034(n27034), .n48(n48), .\read_value[6] (read_value[6]), 
            .n27036(n27036), .n28990(n28990), .\read_value[7] (read_value[7]), 
            .n27028(n27028), .\read_value[8] (read_value[8]), .n27046(n27046), 
            .\read_value[9] (read_value[9]), .n27042(n27042), .\read_value[10] (read_value[10]), 
            .n27045(n27045), .\read_value[11] (read_value[11]), .n27026(n27026), 
            .\read_value[12] (read_value[12]), .n27025(n27025), .\read_value[13] (read_value[13]), 
            .n27027(n27027), .\read_value[14] (read_value[14]), .n27029(n27029), 
            .\read_value[15] (read_value[15]), .n27038(n27038), .\read_value[16] (read_value[16]), 
            .n27031(n27031), .\read_value[17] (read_value[17]), .n27033(n27033), 
            .\read_value[18] (read_value[18]), .n27023(n27023), .\read_value[19] (read_value[19]), 
            .n27041(n27041), .\read_value[20] (read_value[20]), .n27047(n27047), 
            .\read_value[21] (read_value[21]), .n27048(n27048), .\read_value[22] (read_value[22]), 
            .n27040(n27040), .\read_value[23] (read_value[23]), .n27039(n27039), 
            .\read_value[24] (read_value[24]), .n27035(n27035), .\read_value[25] (read_value[25]), 
            .n27050(n27050), .\read_value[26] (read_value[26]), .n27024(n27024), 
            .\read_value[27] (read_value[27]), .n27049(n27049), .\read_value[28] (read_value[28]), 
            .n27044(n27044), .\read_value[29] (read_value[29]), .n27032(n27032), 
            .\read_value[30] (read_value[30]), .n27037(n27037), .\read_value[31] (read_value[31]), 
            .n27043(n27043), .\read_value[0] (read_value[0]), .n14380(n14380), 
            .n27065(n27065), .n14379(n14379), .\databus[1] (databus[1])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(495[45] 505[74])
    LUT4 i1_2_lut_rep_245_3_lut_4_lut (.A(select[4]), .B(n28990), .C(prev_select), 
         .D(n29025), .Z(n28903)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_rep_245_3_lut_4_lut.init = 16'h0002;
    LUT4 Select_3569_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[28]), 
         .D(n30644), .Z(n2)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3569_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i21_2_lut_rep_247_3_lut_4_lut (.A(select[4]), .B(n28990), .C(rw), 
         .D(n26939), .Z(n28905)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i21_2_lut_rep_247_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_3571_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[27]), 
         .D(n30644), .Z(n2_adj_621)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3571_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    VLO i1 (.Z(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i1_4_lut_adj_468 (.A(div_factor_reg_adj_743[8]), .B(n26917), .C(steps_reg_adj_744[8]), 
         .D(register_addr[0]), .Z(n26918)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_468.init = 16'hc088;
    LUT4 Select_3573_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[26]), 
         .D(n30644), .Z(n2_adj_434)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3573_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_260_3_lut_4_lut (.A(select[4]), .B(n28990), .C(prev_select_adj_511), 
         .D(n26939), .Z(n28918)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_rep_260_3_lut_4_lut.init = 16'h0200;
    \ArmPeripheral(axis_haddr=8'b0110000)  arm_a (.databus({databus}), .n3176(n3176), 
            .\register_addr[1] (register_addr[1]), .steps_reg({Open_6, Open_7, 
            Open_8, Open_9, Open_10, Open_11, Open_12, Open_13, 
            Open_14, Open_15, Open_16, Open_17, Open_18, Open_19, 
            Open_20, Open_21, Open_22, Open_23, Open_24, Open_25, 
            Open_26, Open_27, Open_28, Open_29, Open_30, Open_31, 
            Open_32, Open_33, Open_34, Open_35, Open_36, steps_reg_adj_744[0]}), 
            .debug_c_c(debug_c_c), .n30650(n30650), .n15(n15), .\register_addr[0] (register_addr[0]), 
            .VCC_net(VCC_net), .GND_net(GND_net), .Stepper_A_nFault_c(Stepper_A_nFault_c), 
            .\read_size[0] (read_size_adj_746[0]), .n12590(n12590), .n26777(n26777), 
            .n14(n14), .Stepper_A_M0_c_0(Stepper_A_M0_c_0), .n580(n572_adj_684[0]), 
            .\div_factor_reg[0] (div_factor_reg_adj_743[0]), .n12230(n12230), 
            .prev_select(prev_select_adj_551), .n28946(n28946), .n28910(n28910), 
            .n30648(n30648), .n30649(n30649), .\div_factor_reg[4] (div_factor_reg_adj_743[4]), 
            .n609(n581_adj_763[4]), .n611(n581_adj_763[2]), .\control_reg[7] (control_reg_adj_742[7]), 
            .Stepper_A_Dir_c(Stepper_A_Dir_c), .\control_reg[4] (control_reg_adj_742[4]), 
            .Stepper_A_M2_c_2(Stepper_A_M2_c_2), .Stepper_A_M1_c_1(Stepper_A_M1_c_1), 
            .\read_size[2] (read_size_adj_746[2]), .n26870(n26870), .read_value({read_value_adj_745}), 
            .n28929(n28929), .n6120(n6092[4]), .n30651(n30651), .n30652(n30652), 
            .\steps_reg[16] (steps_reg_adj_744[16]), .\steps_reg[8] (steps_reg_adj_744[8]), 
            .\steps_reg[5] (steps_reg_adj_744[5]), .\steps_reg[4] (steps_reg_adj_744[4]), 
            .\steps_reg[3] (steps_reg_adj_744[3]), .n26918(n26918), .stepping(stepping_adj_516), 
            .n30647(n30647), .\div_factor_reg[8] (div_factor_reg_adj_743[8]), 
            .\div_factor_reg[16] (div_factor_reg_adj_743[16]), .n17(n17), 
            .n7(n7), .\select[4] (select[4]), .\register_addr[5] (register_addr[5]), 
            .limit_c_3(limit_c_3), .Stepper_A_En_c(Stepper_A_En_c), .Stepper_A_Step_c(Stepper_A_Step_c), 
            .n24911(n24911), .n26917(n26917), .n27444(n27444), .\register_addr[4] (register_addr[4]), 
            .n11636(n11636), .n28991(n28991)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(604[25] 617[45])
    LUT4 Select_3575_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[25]), 
         .D(n30644), .Z(n2_adj_611)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3575_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i14234_2_lut_2_lut (.A(n30647), .B(databus[0]), .Z(n572_adj_684[0])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14234_2_lut_2_lut.init = 16'h4444;
    LUT4 Select_3577_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[24]), 
         .D(n30644), .Z(n2_adj_624)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3577_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i21240_4_lut (.A(count_adj_802[9]), .B(count_adj_802[11]), .C(count_adj_802[12]), 
         .D(n6_adj_512), .Z(n25126)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i21240_4_lut.init = 16'h0001;
    \ArmPeripheral(axis_haddr=8'b0100000)  arm_z (.read_value({read_value_adj_706}), 
            .debug_c_c(debug_c_c), .n11947(n11947), .GND_net(GND_net), 
            .n30647(n30647), .n28965(n28965), .\register_addr[4] (register_addr[4]), 
            .n28899(n28899), .\register_addr[5] (register_addr[5]), .limit_c_2(limit_c_2), 
            .n7844(n7844), .n14(n14_adj_554), .\register_addr[0] (register_addr[0]), 
            .n15(n15_adj_557), .\register_addr[1] (register_addr[1]), .VCC_net(VCC_net), 
            .Stepper_Z_nFault_c(Stepper_Z_nFault_c), .n30649(n30649), .\read_size[0] (read_size_adj_707[0]), 
            .n84(n84), .Stepper_Z_M0_c_0(Stepper_Z_M0_c_0), .n580(n572_adj_684[0]), 
            .prev_select(prev_select_adj_511), .n28937(n28937), .n30650(n30650), 
            .databus({databus}), .n609(n581_adj_763[4]), .n611(n581_adj_763[2]), 
            .\control_reg[7] (control_reg_adj_703[7]), .n574(n572[6]), .Stepper_Z_Dir_c(Stepper_Z_Dir_c), 
            .Stepper_Z_M2_c_2(Stepper_Z_M2_c_2), .Stepper_Z_M1_c_1(Stepper_Z_M1_c_1), 
            .\read_size[2] (read_size_adj_707[2]), .n60(n60), .n30652(n30652), 
            .n30651(n30651), .\steps_reg[5] (steps_reg_adj_705[5]), .\steps_reg[3] (steps_reg_adj_705[3]), 
            .n29056(n29056), .prev_select_adj_143(prev_select_adj_551), 
            .n28973(n28973), .n12590(n12590), .n29011(n29011), .n29025(n29025), 
            .\register[2][18] (\register[2] [18]), .n29008(n29008), .n27023(n27023), 
            .\register[2][19] (\register[2] [19]), .n27041(n27041), .\register[2][20] (\register[2] [20]), 
            .n27047(n27047), .stepping(stepping_adj_476), .\register[2][21] (\register[2] [21]), 
            .n27048(n27048), .\register[2][22] (\register[2] [22]), .n27040(n27040), 
            .\register[2][23] (\register[2] [23]), .n27039(n27039), .\register[2][24] (\register[2] [24]), 
            .n27035(n27035), .\register[2][25] (\register[2] [25]), .n27050(n27050), 
            .\register[2][26] (\register[2] [26]), .n27024(n27024), .\register[2][27] (\register[2] [27]), 
            .n27049(n27049), .\register[2][28] (\register[2] [28]), .n27044(n27044), 
            .\register[2][29] (\register[2] [29]), .n27032(n27032), .\register[2][30] (\register[2] [30]), 
            .n27037(n27037), .\register[2][31] (\register[2] [31]), .n27043(n27043), 
            .n29021(n29021), .\register_addr[2] (register_addr[2]), .n28955(n28955), 
            .n176(n176), .Stepper_Z_En_c(Stepper_Z_En_c), .Stepper_Z_Step_c(Stepper_Z_Step_c), 
            .rw(rw), .n28956(n28956), .n7(n7), .\register[2][13] (\register[2] [13]), 
            .n27027(n27027), .n30644(n30644), .n28918(n28918), .n26939(n26939), 
            .n27014(n27014), .\register[2][14] (\register[2] [14]), .n27029(n27029), 
            .n24970(n24970), .\register[2][15] (\register[2] [15]), .n27038(n27038), 
            .\register[2][16] (\register[2] [16]), .n27031(n27031), .\register[2][4] (\register[2] [4]), 
            .n27030(n27030), .n28990(n28990), .n11636(n11636), .n26917(n26917), 
            .\register[2][5] (\register[2] [5]), .n27034(n27034), .\register[2][17] (\register[2] [17]), 
            .n27033(n27033), .\register[2][6] (\register[2] [6]), .n27036(n27036), 
            .n22447(n22447), .n27065(n27065), .\register[2][7] (\register[2] [7]), 
            .n27028(n27028), .\register[2][8] (\register[2] [8]), .n27046(n27046), 
            .\register[2][9] (\register[2] [9]), .n27042(n27042), .\register[2][10] (\register[2] [10]), 
            .n27045(n27045), .\register[2][11] (\register[2] [11]), .n27026(n27026), 
            .\register[2][12] (\register[2] [12]), .n27025(n27025), .n28991(n28991)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(589[25] 602[45])
    LUT4 i1_4_lut_adj_469 (.A(register_addr[1]), .B(div_factor_reg_adj_743[16]), 
         .C(steps_reg_adj_744[16]), .D(register_addr[0]), .Z(n17)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_469.init = 16'ha088;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_470 (.A(n30647), .B(prev_select_adj_511), 
         .C(n26939), .D(n28964), .Z(n11947)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_470.init = 16'h1000;
    LUT4 i2_4_lut_4_lut (.A(n30647), .B(n28990), .C(n11618), .D(n28966), 
         .Z(n8050)) /* synthesis lut_function=(!(A+!(B (D)+!B !(C+!(D))))) */ ;
    defparam i2_4_lut_4_lut.init = 16'h4500;
    LUT4 Select_3579_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[23]), 
         .D(n30644), .Z(n2_adj_399)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3579_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i14030_2_lut_2_lut (.A(n30647), .B(n6670), .Z(n241)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14030_2_lut_2_lut.init = 16'h4444;
    LUT4 Select_3581_i2_2_lut_3_lut_4_lut (.A(n28964), .B(n26939), .C(read_value_adj_706[22]), 
         .D(n30644), .Z(n2_adj_626)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3581_i2_2_lut_3_lut_4_lut.init = 16'h8000;
    ClockDivider_U10 pwm_clk_div (.debug_c_c(debug_c_c), .n241(n241), .n30647(n30647), 
            .n6670(n6670), .n27582(n27582), .n24993(n24993), .n28893(n28893), 
            .n27493(n27493), .n24976(n24976), .GND_net(GND_net), .n27569(n27569), 
            .n24988(n24988), .n27575(n27575), .n24998(n24998), .n27590(n27590), 
            .n24991(n24991), .n27548(n27548), .n11996(n11996), .n27556(n27556), 
            .n11997(n11997), .n1018(n1018), .n6(n6_adj_612), .n27509(n27509), 
            .n26690(n26690), .n27527(n27527), .n12104(n12104), .n27640(n27640), 
            .n12804(n12804), .n27638(n27638), .n12807(n12807)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(508[15] 511[41])
    \ArmPeripheral(axis_haddr=8'b0)  arm_x (.\register_addr[1] (register_addr[1]), 
            .\register_addr[0] (register_addr[0]), .databus({databus}), 
            .n3446(n3446), .read_value({read_value_adj_655}), .debug_c_c(debug_c_c), 
            .n11908(n11908), .GND_net(GND_net), .n30651(n30651), .n30648(n30648), 
            .n30649(n30649), .\read_size[0] (read_size_adj_656[0]), .n28920(n28920), 
            .Stepper_X_M0_c_0(Stepper_X_M0_c_0), .n580(n572_adj_684[0]), 
            .prev_select(prev_select), .n28927(n28927), .n30650(n30650), 
            .\steps_reg[7] (steps_reg[7]), .n30652(n30652), .n609(n581_adj_763[4]), 
            .n611(n581_adj_763[2]), .\control_reg[7] (control_reg[7]), .n574(n572[6]), 
            .Stepper_X_Dir_c(Stepper_X_Dir_c), .Stepper_X_M2_c_2(Stepper_X_M2_c_2), 
            .Stepper_X_M1_c_1(Stepper_X_M1_c_1), .\read_size[2] (read_size_adj_656[2]), 
            .n28901(n28901), .n30653(n30653), .n28991(n28991), .rw(rw), 
            .n28903(n28903), .n29052(n29052), .n28917(n28917), .Stepper_X_En_c(Stepper_X_En_c), 
            .Stepper_X_Step_c(Stepper_X_Step_c), .limit_c_0(limit_c_0), 
            .n29025(n29025), .n30647(n30647), .n28898(n28898), .n28965(n28965), 
            .n24994(n24994), .n21(n21), .VCC_net(VCC_net), .Stepper_X_nFault_c(Stepper_X_nFault_c), 
            .n13(n13)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(559[25] 572[45])
    RCPeripheral rc_receiver (.databus_out({databus_out}), .n2(n2_adj_585), 
            .rw(rw), .databus({databus}), .\read_value[9] (read_value[9]), 
            .n1(n1_adj_584), .n29028(n29028), .\read_value[9]_adj_1 (read_value_adj_655[9]), 
            .read_value({read_value_adj_667}), .n28904(n28904), .n53(n53), 
            .n2_adj_3(n2_adj_581), .\read_value[8]_adj_4 (read_value[8]), 
            .n1_adj_5(n1_adj_580), .\read_value[8]_adj_6 (read_value_adj_655[8]), 
            .\register_addr[0] (register_addr[0]), .n4(n4_adj_587), .\read_value[7]_adj_7 (read_value_adj_745[7]), 
            .n28928(n28928), .\select[7] (select[7]), .\read_value[7]_adj_8 (read_value_adj_706[7]), 
            .\read_value[7]_adj_9 (read_value[7]), .n28905(n28905), .n30644(n30644), 
            .read_value_adj_142({read_value_adj_650}), .n64(n64), .n4_adj_18(n4_adj_586), 
            .n176(n176), .\read_value[6]_adj_19 (read_value_adj_745[6]), 
            .\read_value[6]_adj_20 (read_value_adj_706[6]), .\read_value[6]_adj_21 (read_value[6]), 
            .n2_adj_22(n2_adj_597), .\read_value[17]_adj_23 (read_value[17]), 
            .n1_adj_24(n1_adj_596), .\read_value[17]_adj_25 (read_value_adj_655[17]), 
            .n2_adj_26(n2_adj_605), .\read_value[16]_adj_27 (read_value[16]), 
            .n1_adj_28(n1_adj_604), .\read_value[16]_adj_29 (read_value_adj_655[16]), 
            .n2_adj_30(n2_adj_603), .\read_value[15]_adj_31 (read_value[15]), 
            .n1_adj_32(n1_adj_602), .\read_value[15]_adj_33 (read_value_adj_655[15]), 
            .n2_adj_34(n2_adj_593), .\read_value[14]_adj_35 (read_value[14]), 
            .n1_adj_36(n1_adj_592), .\read_value[14]_adj_37 (read_value_adj_655[14]), 
            .n4_adj_38(n4_adj_577), .\read_value[5]_adj_39 (read_value_adj_745[5]), 
            .\read_value[5]_adj_40 (read_value_adj_706[5]), .\read_value[5]_adj_41 (read_value[5]), 
            .n2_adj_42(n2_adj_591), .\read_value[13]_adj_43 (read_value[13]), 
            .n1_adj_44(n1_adj_590), .\register_addr[2] (register_addr[2]), 
            .\read_value[13]_adj_45 (read_value_adj_655[13]), .n2_adj_46(n2_adj_561), 
            .\read_value[31]_adj_47 (read_value[31]), .n1_adj_48(n1_adj_562), 
            .\read_value[31]_adj_49 (read_value_adj_655[31]), .n2_adj_50(n2_adj_627), 
            .\read_value[30]_adj_51 (read_value[30]), .n1_adj_52(n1_adj_472), 
            .n2_adj_53(n2_adj_589), .\read_value[12]_adj_54 (read_value[12]), 
            .n1_adj_55(n1_adj_588), .\read_value[12]_adj_56 (read_value_adj_655[12]), 
            .\read_value[30]_adj_57 (read_value_adj_655[30]), .\register_addr[1] (register_addr[1]), 
            .n2_adj_58(n2_adj_608), .\read_value[29]_adj_59 (read_value[29]), 
            .n1_adj_60(n1_adj_552), .\read_value[29]_adj_61 (read_value_adj_655[29]), 
            .n2_adj_62(n2_adj_583), .\read_value[11]_adj_63 (read_value[11]), 
            .n1_adj_64(n1_adj_582), .\read_value[11]_adj_65 (read_value_adj_655[11]), 
            .n2_adj_66(n2_adj_579), .\read_value[10]_adj_67 (read_value[10]), 
            .n1_adj_68(n1_adj_578), .\read_value[10]_adj_69 (read_value_adj_655[10]), 
            .n28955(n28955), .read_size({read_size}), .\select[1] (select[1]), 
            .n29018(n29018), .\sendcount[1] (sendcount[1]), .n11253(n11253), 
            .\read_size[2]_adj_70 (read_size_adj_707[2]), .n28937(n28937), 
            .\reg_size[2] (reg_size[2]), .n28946(n28946), .\read_size[2]_adj_71 (read_size_adj_746[2]), 
            .n4_adj_72(n4_adj_576), .\read_value[4]_adj_73 (read_value_adj_745[4]), 
            .\read_value[4]_adj_74 (read_value_adj_706[4]), .\read_value[4]_adj_75 (read_value[4]), 
            .n2_adj_76(n2), .\read_value[28]_adj_77 (read_value[28]), .n1_adj_78(n1_adj_471), 
            .\read_value[28]_adj_79 (read_value_adj_655[28]), .n2_adj_80(n2_adj_621), 
            .\read_value[27]_adj_81 (read_value[27]), .n1_adj_82(n1_adj_389), 
            .\read_value[27]_adj_83 (read_value_adj_655[27]), .n2_adj_84(n2_adj_434), 
            .n4_adj_85(n4_adj_565), .\read_value[26]_adj_86 (read_value[26]), 
            .n1_adj_87(n1_adj_390), .\read_value[3]_adj_88 (read_value_adj_745[3]), 
            .\read_value[26]_adj_89 (read_value_adj_655[26]), .n2_adj_90(n2_adj_611), 
            .\read_value[3]_adj_91 (read_value_adj_706[3]), .\read_value[3]_adj_92 (read_value[3]), 
            .\read_value[25]_adj_93 (read_value[25]), .n1_adj_94(n1_adj_553), 
            .\read_value[25]_adj_95 (read_value_adj_655[25]), .n2_adj_96(n2_adj_624), 
            .\read_value[24]_adj_97 (read_value[24]), .n1_adj_98(n1_adj_623), 
            .\read_value[24]_adj_99 (read_value_adj_655[24]), .n4_adj_100(n4_adj_564), 
            .\read_value[2]_adj_101 (read_value_adj_745[2]), .n2_adj_102(n2_adj_399), 
            .\read_value[2]_adj_103 (read_value_adj_706[2]), .\read_value[2]_adj_104 (read_value[2]), 
            .\read_value[23]_adj_105 (read_value[23]), .n1_adj_106(n1_adj_625), 
            .\read_value[23]_adj_107 (read_value_adj_655[23]), .n2_adj_108(n2_adj_626), 
            .n1_adj_109(n1_adj_566), .\read_value[22]_adj_110 (read_value[22]), 
            .n1_adj_111(n1), .\read_value[1]_adj_112 (read_value_adj_655[1]), 
            .n6(n6_adj_567), .\read_value[22]_adj_113 (read_value_adj_655[22]), 
            .n2_adj_114(n2_adj_607), .\read_value[1]_adj_115 (read_value_adj_706[1]), 
            .\read_value[21]_adj_116 (read_value[21]), .n1_adj_117(n1_adj_606), 
            .\read_value[21]_adj_118 (read_value_adj_655[21]), .n2_adj_119(n2_adj_599), 
            .\read_value[20]_adj_120 (read_value[20]), .n1_adj_121(n1_adj_598), 
            .\read_value[20]_adj_122 (read_value_adj_655[20]), .n4_adj_123(n4_adj_563), 
            .\read_value[0]_adj_124 (read_value_adj_745[0]), .\read_value[0]_adj_125 (read_value_adj_706[0]), 
            .\read_value[0]_adj_126 (read_value[0]), .\read_size[2]_adj_127 (read_size_adj_656[2]), 
            .\read_size[2]_adj_128 (read_size_adj_668[2]), .n28927(n28927), 
            .n28974(n28974), .\read_size[0]_adj_129 (read_size_adj_707[0]), 
            .n9(n9), .\read_size[0]_adj_130 (read_size_adj_668[0]), .\read_size[0]_adj_131 (read_size_adj_746[0]), 
            .n10(n10_adj_560), .\read_size[0]_adj_132 (read_size_adj_651[0]), 
            .\select[2] (select[2]), .n8(n8), .n2_adj_133(n2_adj_595), 
            .\read_value[19]_adj_134 (read_value[19]), .n1_adj_135(n1_adj_594), 
            .n2_adj_136(n2_adj_601), .\read_value[19]_adj_137 (read_value_adj_655[19]), 
            .\read_value[18]_adj_138 (read_value[18]), .n1_adj_139(n1_adj_600), 
            .\read_value[18]_adj_140 (read_value_adj_655[18]), .debug_c_c(debug_c_c), 
            .n28893(n28893), .rc_ch8_c(rc_ch8_c), .GND_net(GND_net), .n27548(n27548), 
            .n27590(n27590), .n11996(n11996), .n24991(n24991), .n27575(n27575), 
            .rc_ch7_c(rc_ch7_c), .n11997(n11997), .n27556(n27556), .n24998(n24998), 
            .n1030(n1030), .n1018(n1018), .n27509(n27509), .n4_adj_141(n4_adj_558), 
            .rc_ch4_c(rc_ch4_c), .n54(n54), .n26690(n26690), .n28888(n28888), 
            .n14053(n14053), .n27569(n27569), .rc_ch3_c(rc_ch3_c), .n27527(n27527), 
            .n12104(n12104), .n24988(n24988), .n27582(n27582), .n27640(n27640), 
            .n12804(n12804), .rc_ch2_c(rc_ch2_c), .n24993(n24993), .n27493(n27493), 
            .n27638(n27638), .n12807(n12807), .rc_ch1_c(rc_ch1_c), .n24976(n24976)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(622[15] 634[41])
    
endmodule
//
// Verilog Description of module PWMPeripheral
//

module PWMPeripheral (\read_size[0] , debug_c_c, n28920, n30649, \databus[0] , 
            \select[2] , n282, n30653, \databus[6] , \databus[5] , 
            \databus[4] , \databus[3] , \databus[2] , \databus[1] , 
            n29063, n28900, n30647, \register_addr[0] , rw, read_value, 
            n8044, n64, \count[0] , n10489, n28893, GND_net, n7885, 
            n7894, \count[3] , n14286, \count[7] , \count[5] , \count[1] , 
            \count[6] , \count[8] , \count[4] , \count[2] , motor_pwm_r_c, 
            n3585, \count[0]_adj_185 , n10501, n14439, \count[12] , 
            \count[11] , \count[9] , \count[8]_adj_186 , \count[6]_adj_187 , 
            \count[5]_adj_188 , \count[3]_adj_189 , \count[2]_adj_190 , 
            \count[1]_adj_191 , n28911, n10, n12, \reset_count[5] , 
            n27079, \reset_count[6] , \reset_count[4] , n27080, \reset_count[8] , 
            \reset_count[7] , n7904, n7898, n7897, n7900, n7902, 
            n7901, n7903, motor_pwm_l_c, n25126, n28958, n6, n8, 
            n3582, n6_adj_192) /* synthesis syn_module_defined=1 */ ;
    output \read_size[0] ;
    input debug_c_c;
    input n28920;
    input n30649;
    input \databus[0] ;
    input \select[2] ;
    input n282;
    input n30653;
    input \databus[6] ;
    input \databus[5] ;
    input \databus[4] ;
    input \databus[3] ;
    input \databus[2] ;
    input \databus[1] ;
    output n29063;
    input n28900;
    input n30647;
    input \register_addr[0] ;
    input rw;
    output [7:0]read_value;
    input n8044;
    output n64;
    output \count[0] ;
    output n10489;
    input n28893;
    input GND_net;
    output [7:0]n7885;
    output n7894;
    output \count[3] ;
    input n14286;
    output \count[7] ;
    output \count[5] ;
    output \count[1] ;
    output \count[6] ;
    output \count[8] ;
    output \count[4] ;
    output \count[2] ;
    output motor_pwm_r_c;
    input n3585;
    output \count[0]_adj_185 ;
    output n10501;
    input n14439;
    output \count[12] ;
    output \count[11] ;
    output \count[9] ;
    output \count[8]_adj_186 ;
    output \count[6]_adj_187 ;
    output \count[5]_adj_188 ;
    output \count[3]_adj_189 ;
    output \count[2]_adj_190 ;
    output \count[1]_adj_191 ;
    output n28911;
    input n10;
    output n12;
    input \reset_count[5] ;
    output n27079;
    input \reset_count[6] ;
    input \reset_count[4] ;
    output n27080;
    input \reset_count[8] ;
    input \reset_count[7] ;
    output n7904;
    output n7898;
    output n7897;
    output n7900;
    output n7902;
    output n7901;
    output n7903;
    output motor_pwm_l_c;
    input n25126;
    output n28958;
    input n6;
    output n8;
    input n3582;
    output n6_adj_192;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n12065;
    wire [7:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(55[12:20])
    
    wire n28895, prev_select;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(55[12:20])
    
    wire n12532, n28894, n20619;
    wire [7:0]n4890;
    
    FD1P3AX read_size__i1 (.D(n28920), .SP(n12065), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3JX register_0__i1 (.D(\databus[0] ), .SP(n28895), .PD(n30649), 
            .CK(debug_c_c), .Q(\register[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i1.GSR = "ENABLED";
    FD1S3AX prev_select_138 (.D(\select[2] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam prev_select_138.GSR = "ENABLED";
    FD1P3AX register_0__i16 (.D(n282), .SP(n12532), .CK(debug_c_c), .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i16.GSR = "ENABLED";
    FD1P3JX register_0__i15 (.D(\databus[6] ), .SP(n28894), .PD(n30653), 
            .CK(debug_c_c), .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i15.GSR = "ENABLED";
    FD1P3JX register_0__i14 (.D(\databus[5] ), .SP(n28894), .PD(n30653), 
            .CK(debug_c_c), .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i14.GSR = "ENABLED";
    FD1P3JX register_0__i13 (.D(\databus[4] ), .SP(n28894), .PD(n30653), 
            .CK(debug_c_c), .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i13.GSR = "ENABLED";
    FD1P3JX register_0__i12 (.D(\databus[3] ), .SP(n28894), .PD(n30653), 
            .CK(debug_c_c), .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i12.GSR = "ENABLED";
    FD1P3JX register_0__i11 (.D(\databus[2] ), .SP(n28894), .PD(n30653), 
            .CK(debug_c_c), .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i11.GSR = "ENABLED";
    FD1P3JX register_0__i10 (.D(\databus[1] ), .SP(n28894), .PD(n30653), 
            .CK(debug_c_c), .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i10.GSR = "ENABLED";
    FD1P3JX register_0__i9 (.D(\databus[0] ), .SP(n28894), .PD(n30653), 
            .CK(debug_c_c), .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i9.GSR = "ENABLED";
    FD1P3AX register_0__i8 (.D(n282), .SP(n20619), .CK(debug_c_c), .Q(\register[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i8.GSR = "ENABLED";
    FD1P3JX register_0__i7 (.D(\databus[6] ), .SP(n28895), .PD(n30653), 
            .CK(debug_c_c), .Q(\register[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i7.GSR = "ENABLED";
    FD1P3JX register_0__i6 (.D(\databus[5] ), .SP(n28895), .PD(n30653), 
            .CK(debug_c_c), .Q(\register[0] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i6.GSR = "ENABLED";
    FD1P3JX register_0__i5 (.D(\databus[4] ), .SP(n28895), .PD(n30653), 
            .CK(debug_c_c), .Q(\register[0] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i5.GSR = "ENABLED";
    FD1P3JX register_0__i4 (.D(\databus[3] ), .SP(n28895), .PD(n30653), 
            .CK(debug_c_c), .Q(\register[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i4.GSR = "ENABLED";
    FD1P3JX register_0__i3 (.D(\databus[2] ), .SP(n28895), .PD(n30653), 
            .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i3.GSR = "ENABLED";
    FD1P3JX register_0__i2 (.D(\databus[1] ), .SP(n28895), .PD(n30653), 
            .CK(debug_c_c), .Q(\register[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i2.GSR = "ENABLED";
    LUT4 i21243_2_lut_3_lut_4_lut (.A(n29063), .B(n28900), .C(n30647), 
         .D(\register_addr[0] ), .Z(n20619)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C)) */ ;
    defparam i21243_2_lut_3_lut_4_lut.init = 16'hf0f2;
    LUT4 i1_2_lut_rep_405 (.A(\select[2] ), .B(prev_select), .Z(n29063)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(82[8:29])
    defparam i1_2_lut_rep_405.init = 16'h2222;
    LUT4 i1_2_lut_2_lut_3_lut (.A(\select[2] ), .B(prev_select), .C(n30647), 
         .Z(n12065)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(82[8:29])
    defparam i1_2_lut_2_lut_3_lut.init = 16'h0202;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n29063), .B(n28900), .C(n30647), .D(\register_addr[0] ), 
         .Z(n12532)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf2f0;
    LUT4 i3864_2_lut_rep_236_3_lut_4_lut (.A(rw), .B(n28920), .C(\register_addr[0] ), 
         .D(n29063), .Z(n28894)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i3864_2_lut_rep_236_3_lut_4_lut.init = 16'h4000;
    LUT4 i21251_2_lut_rep_237_3_lut_4_lut (.A(rw), .B(n28920), .C(\register_addr[0] ), 
         .D(n29063), .Z(n28895)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i21251_2_lut_rep_237_3_lut_4_lut.init = 16'h0400;
    FD1P3IX read_value__i0 (.D(n4890[0]), .SP(n12065), .CD(n8044), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 mux_1582_Mux_0_i1_3_lut (.A(\register[0] [0]), .B(\register[1] [0]), 
         .C(\register_addr[0] ), .Z(n4890[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1582_Mux_0_i1_3_lut.init = 16'hcaca;
    LUT4 i16_2_lut (.A(\select[2] ), .B(rw), .Z(n64)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(68[19:32])
    defparam i16_2_lut.init = 16'h8888;
    LUT4 mux_1582_Mux_1_i1_3_lut (.A(\register[0] [1]), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n4890[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1582_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1582_Mux_2_i1_3_lut (.A(\register[0] [2]), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n4890[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1582_Mux_2_i1_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i1 (.D(n4890[1]), .SP(n12065), .CD(n8044), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n4890[2]), .SP(n12065), .CD(n8044), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n4890[3]), .SP(n12065), .CD(n8044), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n4890[4]), .SP(n12065), .CD(n8044), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n4890[5]), .SP(n12065), .CD(n8044), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n4890[6]), .SP(n12065), .CD(n8044), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n4890[7]), .SP(n12065), .CD(n8044), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i7.GSR = "ENABLED";
    LUT4 mux_1582_Mux_3_i1_3_lut (.A(\register[0] [3]), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n4890[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1582_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1582_Mux_4_i1_3_lut (.A(\register[0] [4]), .B(\register[1] [4]), 
         .C(\register_addr[0] ), .Z(n4890[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1582_Mux_4_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1582_Mux_5_i1_3_lut (.A(\register[0] [5]), .B(\register[1] [5]), 
         .C(\register_addr[0] ), .Z(n4890[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1582_Mux_5_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1582_Mux_6_i1_3_lut (.A(\register[0] [6]), .B(\register[1] [6]), 
         .C(\register_addr[0] ), .Z(n4890[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1582_Mux_6_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1582_Mux_7_i1_3_lut (.A(\register[0] [7]), .B(\register[1] [7]), 
         .C(\register_addr[0] ), .Z(n4890[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1582_Mux_7_i1_3_lut.init = 16'hcaca;
    PWMGenerator right (.count({Open_37, Open_38, Open_39, Open_40, 
            Open_41, Open_42, Open_43, Open_44, Open_45, Open_46, 
            Open_47, Open_48, \count[0] }), .n10489(n10489), .n28893(n28893), 
            .debug_c_c(debug_c_c), .GND_net(GND_net), .n7885({n7885}), 
            .n7894(n7894), .\count[3] (\count[3] ), .n14286(n14286), .\register[1] ({\register[1] }), 
            .n30647(n30647), .\count[7] (\count[7] ), .\count[5] (\count[5] ), 
            .\count[1] (\count[1] ), .\count[6] (\count[6] ), .\count[8] (\count[8] ), 
            .\count[4] (\count[4] ), .\count[2] (\count[2] ), .motor_pwm_r_c(motor_pwm_r_c), 
            .n3585(n3585)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(118[15] 121[34])
    PWMGenerator_U6 left (.count({\count[12] , \count[11] , Open_49, Open_50, 
            Open_51, Open_52, Open_53, Open_54, Open_55, Open_56, 
            Open_57, Open_58, \count[0]_adj_185 }), .debug_c_c(debug_c_c), 
            .n28893(n28893), .n10501(n10501), .n14439(n14439), .\register[0] ({\register[0] }), 
            .\count[9] (\count[9] ), .\count[8] (\count[8]_adj_186 ), .\count[6] (\count[6]_adj_187 ), 
            .\count[5] (\count[5]_adj_188 ), .\count[3] (\count[3]_adj_189 ), 
            .\count[2] (\count[2]_adj_190 ), .\count[1] (\count[1]_adj_191 ), 
            .n28911(n28911), .n10(n10), .n12(n12), .\reset_count[5] (\reset_count[5] ), 
            .n27079(n27079), .\reset_count[6] (\reset_count[6] ), .\reset_count[4] (\reset_count[4] ), 
            .n27080(n27080), .\reset_count[8] (\reset_count[8] ), .\reset_count[7] (\reset_count[7] ), 
            .n30647(n30647), .GND_net(GND_net), .n7904(n7904), .n7898(n7898), 
            .n7897(n7897), .n7900(n7900), .n7902(n7902), .n7901(n7901), 
            .n7903(n7903), .motor_pwm_l_c(motor_pwm_l_c), .n25126(n25126), 
            .n28958(n28958), .n6(n6), .n8(n8), .n3582(n3582), .n6_adj_184(n6_adj_192)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(114[15] 117[34])
    
endmodule
//
// Verilog Description of module PWMGenerator
//

module PWMGenerator (count, n10489, n28893, debug_c_c, GND_net, n7885, 
            n7894, \count[3] , n14286, \register[1] , n30647, \count[7] , 
            \count[5] , \count[1] , \count[6] , \count[8] , \count[4] , 
            \count[2] , motor_pwm_r_c, n3585) /* synthesis syn_module_defined=1 */ ;
    output [12:0]count;
    output n10489;
    input n28893;
    input debug_c_c;
    input GND_net;
    output [7:0]n7885;
    output n7894;
    output \count[3] ;
    input n14286;
    input [7:0]\register[1] ;
    input n30647;
    output \count[7] ;
    output \count[5] ;
    output \count[1] ;
    output \count[6] ;
    output \count[8] ;
    output \count[4] ;
    output \count[2] ;
    output motor_pwm_r_c;
    input n3585;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n7, n27197, n20039, n27273, n27337, n27287, n8023;
    wire [12:0]n43;
    
    wire n24252;
    wire [7:0]latched_width;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(15[12:25])
    
    wire n24251;
    wire [12:0]count_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    
    wire n24250, n24249, n26897, n17, n16;
    wire [12:0]n28;
    
    wire n24588, n24587, n24586, n24585, n24584, n24583, n25181;
    
    LUT4 i4_4_lut (.A(n7), .B(n27197), .C(n20039), .D(count[0]), .Z(n10489)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i4_4_lut.init = 16'h0002;
    LUT4 i2_4_lut (.A(n27273), .B(n28893), .C(n27337), .D(n27287), .Z(n7)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i2_4_lut.init = 16'h0004;
    FD1P3IX count__i0 (.D(n43[0]), .SP(n28893), .CD(n8023), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i0.GSR = "ENABLED";
    CCU2D add_2153_9 (.A0(latched_width[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24252), .S0(n7885[7]), .S1(n7894));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2153_9.INIT0 = 16'h5555;
    defparam add_2153_9.INIT1 = 16'h0000;
    defparam add_2153_9.INJECT1_0 = "NO";
    defparam add_2153_9.INJECT1_1 = "NO";
    CCU2D add_2153_7 (.A0(latched_width[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24251), .COUT(n24252), .S0(n7885[5]), 
          .S1(n7885[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2153_7.INIT0 = 16'h5555;
    defparam add_2153_7.INIT1 = 16'h5555;
    defparam add_2153_7.INJECT1_0 = "NO";
    defparam add_2153_7.INJECT1_1 = "NO";
    LUT4 i20903_2_lut (.A(count_c[9]), .B(\count[3] ), .Z(n27273)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20903_2_lut.init = 16'heeee;
    FD1P3JX latched_width_i0_i2 (.D(\register[1] [2]), .SP(n10489), .PD(n14286), 
            .CK(debug_c_c), .Q(latched_width[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i2.GSR = "ENABLED";
    CCU2D add_2153_5 (.A0(latched_width[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24250), .COUT(n24251), .S0(n7885[3]), 
          .S1(n7885[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2153_5.INIT0 = 16'h5555;
    defparam add_2153_5.INIT1 = 16'h5555;
    defparam add_2153_5.INJECT1_0 = "NO";
    defparam add_2153_5.INJECT1_1 = "NO";
    CCU2D add_2153_3 (.A0(latched_width[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24249), .COUT(n24250), .S0(n7885[1]), 
          .S1(n7885[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2153_3.INIT0 = 16'h5555;
    defparam add_2153_3.INIT1 = 16'h5555;
    defparam add_2153_3.INJECT1_0 = "NO";
    defparam add_2153_3.INJECT1_1 = "NO";
    LUT4 i2266_4_lut (.A(n28893), .B(n26897), .C(n30647), .D(n20039), 
         .Z(n8023)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam i2266_4_lut.init = 16'ha0a8;
    FD1P3JX latched_width_i0_i3 (.D(\register[1] [3]), .SP(n10489), .PD(n14286), 
            .CK(debug_c_c), .Q(latched_width[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i3.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i4 (.D(\register[1] [4]), .SP(n10489), .PD(n14286), 
            .CK(debug_c_c), .Q(latched_width[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i4.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i5 (.D(\register[1] [5]), .SP(n10489), .PD(n14286), 
            .CK(debug_c_c), .Q(latched_width[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i5.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i6 (.D(\register[1] [6]), .SP(n10489), .PD(n14286), 
            .CK(debug_c_c), .Q(latched_width[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i6.GSR = "ENABLED";
    LUT4 i20967_4_lut (.A(\count[7] ), .B(\count[5] ), .C(\count[1] ), 
         .D(count_c[12]), .Z(n27337)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20967_4_lut.init = 16'hfffe;
    LUT4 i20917_2_lut (.A(\count[6] ), .B(\count[8] ), .Z(n27287)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20917_2_lut.init = 16'heeee;
    CCU2D add_2153_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(latched_width[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24249), .S1(n7885[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2153_1.INIT0 = 16'hF000;
    defparam add_2153_1.INIT1 = 16'h5555;
    defparam add_2153_1.INJECT1_0 = "NO";
    defparam add_2153_1.INJECT1_1 = "NO";
    LUT4 i9_4_lut (.A(n17), .B(\count[5] ), .C(n16), .D(n27197), .Z(n26897)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i9_4_lut.init = 16'h0080;
    LUT4 i7_4_lut (.A(count[0]), .B(count_c[9]), .C(count_c[12]), .D(\count[6] ), 
         .Z(n17)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(\count[7] ), .B(\count[8] ), .C(\count[3] ), .D(\count[1] ), 
         .Z(n16)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i20833_2_lut (.A(count_c[10]), .B(count_c[11]), .Z(n27197)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20833_2_lut.init = 16'heeee;
    FD1P3IX count__i11 (.D(n28[11]), .SP(n28893), .CD(n8023), .CK(debug_c_c), 
            .Q(count_c[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n28[12]), .SP(n28893), .CD(n8023), .CK(debug_c_c), 
            .Q(count_c[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i12.GSR = "ENABLED";
    LUT4 i14309_2_lut (.A(\count[4] ), .B(\count[2] ), .Z(n20039)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14309_2_lut.init = 16'heeee;
    CCU2D add_9_13 (.A0(count_c[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24588), .S0(n28[11]), .S1(n28[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_13.INIT0 = 16'h5aaa;
    defparam add_9_13.INIT1 = 16'h5aaa;
    defparam add_9_13.INJECT1_0 = "NO";
    defparam add_9_13.INJECT1_1 = "NO";
    CCU2D add_9_11 (.A0(count_c[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24587), .COUT(n24588), .S0(n28[9]), .S1(n28[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_11.INIT0 = 16'h5aaa;
    defparam add_9_11.INIT1 = 16'h5aaa;
    defparam add_9_11.INJECT1_0 = "NO";
    defparam add_9_11.INJECT1_1 = "NO";
    CCU2D add_9_9 (.A0(\count[7] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count[8] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24586), .COUT(n24587), .S0(n28[7]), .S1(n28[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_9.INIT0 = 16'h5aaa;
    defparam add_9_9.INIT1 = 16'h5aaa;
    defparam add_9_9.INJECT1_0 = "NO";
    defparam add_9_9.INJECT1_1 = "NO";
    FD1P3IX latched_width_i0_i7 (.D(\register[1] [7]), .SP(n10489), .CD(n14286), 
            .CK(debug_c_c), .Q(latched_width[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i7.GSR = "ENABLED";
    CCU2D add_9_7 (.A0(\count[5] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count[6] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24585), .COUT(n24586), .S0(n28[5]), .S1(n28[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_7.INIT0 = 16'h5aaa;
    defparam add_9_7.INIT1 = 16'h5aaa;
    defparam add_9_7.INJECT1_0 = "NO";
    defparam add_9_7.INJECT1_1 = "NO";
    CCU2D add_9_5 (.A0(\count[3] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count[4] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24584), .COUT(n24585), .S0(n28[3]), .S1(n28[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_5.INIT0 = 16'h5aaa;
    defparam add_9_5.INIT1 = 16'h5aaa;
    defparam add_9_5.INJECT1_0 = "NO";
    defparam add_9_5.INJECT1_1 = "NO";
    CCU2D add_9_3 (.A0(\count[1] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count[2] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24583), .COUT(n24584), .S0(n28[1]), .S1(n28[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_3.INIT0 = 16'h5aaa;
    defparam add_9_3.INIT1 = 16'h5aaa;
    defparam add_9_3.INJECT1_0 = "NO";
    defparam add_9_3.INJECT1_1 = "NO";
    CCU2D add_9_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24583), 
          .S1(n43[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_1.INIT0 = 16'hF000;
    defparam add_9_1.INIT1 = 16'h5555;
    defparam add_9_1.INJECT1_0 = "NO";
    defparam add_9_1.INJECT1_1 = "NO";
    OFS1P3IX pwm_19 (.D(n25181), .SP(n28893), .SCLK(debug_c_c), .CD(GND_net), 
            .Q(motor_pwm_r_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam pwm_19.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i0 (.D(\register[1] [0]), .SP(n10489), .PD(n14286), 
            .CK(debug_c_c), .Q(latched_width[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i0.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i1 (.D(\register[1] [1]), .SP(n10489), .PD(n14286), 
            .CK(debug_c_c), .Q(latched_width[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i1.GSR = "ENABLED";
    LUT4 i21342_4_lut (.A(n27197), .B(count_c[12]), .C(n3585), .D(count_c[9]), 
         .Z(n25181)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(31[7:16])
    defparam i21342_4_lut.init = 16'h0001;
    FD1P3IX count__i1 (.D(n28[1]), .SP(n28893), .CD(n8023), .CK(debug_c_c), 
            .Q(\count[1] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i1.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n28[2]), .SP(n28893), .CD(n8023), .CK(debug_c_c), 
            .Q(\count[2] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n28[3]), .SP(n28893), .CD(n8023), .CK(debug_c_c), 
            .Q(\count[3] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n28[4]), .SP(n28893), .CD(n8023), .CK(debug_c_c), 
            .Q(\count[4] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n28[5]), .SP(n28893), .CD(n8023), .CK(debug_c_c), 
            .Q(\count[5] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n28[6]), .SP(n28893), .CD(n8023), .CK(debug_c_c), 
            .Q(\count[6] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n28[7]), .SP(n28893), .CD(n8023), .CK(debug_c_c), 
            .Q(\count[7] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n28[8]), .SP(n28893), .CD(n8023), .CK(debug_c_c), 
            .Q(\count[8] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n28[9]), .SP(n28893), .CD(n8023), .CK(debug_c_c), 
            .Q(count_c[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n28[10]), .SP(n28893), .CD(n8023), .CK(debug_c_c), 
            .Q(count_c[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i10.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMGenerator_U6
//

module PWMGenerator_U6 (count, debug_c_c, n28893, n10501, n14439, 
            \register[0] , \count[9] , \count[8] , \count[6] , \count[5] , 
            \count[3] , \count[2] , \count[1] , n28911, n10, n12, 
            \reset_count[5] , n27079, \reset_count[6] , \reset_count[4] , 
            n27080, \reset_count[8] , \reset_count[7] , n30647, GND_net, 
            n7904, n7898, n7897, n7900, n7902, n7901, n7903, motor_pwm_l_c, 
            n25126, n28958, n6, n8, n3582, n6_adj_184) /* synthesis syn_module_defined=1 */ ;
    output [12:0]count;
    input debug_c_c;
    input n28893;
    output n10501;
    input n14439;
    input [7:0]\register[0] ;
    output \count[9] ;
    output \count[8] ;
    output \count[6] ;
    output \count[5] ;
    output \count[3] ;
    output \count[2] ;
    output \count[1] ;
    output n28911;
    input n10;
    output n12;
    input \reset_count[5] ;
    output n27079;
    input \reset_count[6] ;
    input \reset_count[4] ;
    output n27080;
    input \reset_count[8] ;
    input \reset_count[7] ;
    input n30647;
    input GND_net;
    output n7904;
    output n7898;
    output n7897;
    output n7900;
    output n7902;
    output n7901;
    output n7903;
    output motor_pwm_l_c;
    input n25126;
    output n28958;
    input n6;
    output n8;
    input n3582;
    output n6_adj_184;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [12:0]n42;
    wire [7:0]latched_width;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(15[12:25])
    
    wire n8019;
    wire [12:0]n43;
    wire [12:0]count_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    
    wire n27223, n20;
    wire [7:0]n7895;
    wire [12:0]n28;
    
    wire n25195, n15_adj_378, n14, n27347, n27327, n27231, n24581, 
        n24580, n24579, n24578, n24577, n24576, n24575, n24574, 
        n24573, n24572;
    
    FD1P3AX count__i0 (.D(n42[0]), .SP(n28893), .CK(debug_c_c), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i0.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i0 (.D(\register[0] [0]), .SP(n10501), .PD(n14439), 
            .CK(debug_c_c), .Q(latched_width[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i0.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n43[12]), .SP(n28893), .CD(n8019), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i12.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n43[11]), .SP(n28893), .CD(n8019), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n43[10]), .SP(n28893), .CD(n8019), .CK(debug_c_c), 
            .Q(count_c[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n43[9]), .SP(n28893), .CD(n8019), .CK(debug_c_c), 
            .Q(\count[9] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n43[8]), .SP(n28893), .CD(n8019), .CK(debug_c_c), 
            .Q(\count[8] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n43[7]), .SP(n28893), .CD(n8019), .CK(debug_c_c), 
            .Q(count_c[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n43[6]), .SP(n28893), .CD(n8019), .CK(debug_c_c), 
            .Q(\count[6] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n43[5]), .SP(n28893), .CD(n8019), .CK(debug_c_c), 
            .Q(\count[5] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n43[4]), .SP(n28893), .CD(n8019), .CK(debug_c_c), 
            .Q(count_c[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n43[3]), .SP(n28893), .CD(n8019), .CK(debug_c_c), 
            .Q(\count[3] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n43[2]), .SP(n28893), .CD(n8019), .CK(debug_c_c), 
            .Q(\count[2] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n43[1]), .SP(n28893), .CD(n8019), .CK(debug_c_c), 
            .Q(\count[1] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i1.GSR = "ENABLED";
    LUT4 i20857_3_lut_4_lut (.A(\count[2] ), .B(count_c[4]), .C(count[11]), 
         .D(count_c[10]), .Z(n27223)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20857_3_lut_4_lut.init = 16'hfffe;
    LUT4 i7_3_lut_4_lut (.A(\count[2] ), .B(count_c[4]), .C(\count[8] ), 
         .D(n28893), .Z(n20)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i7_3_lut_4_lut.init = 16'h0100;
    LUT4 i10_2_lut_rep_253 (.A(n7895[7]), .B(count_c[7]), .Z(n28911)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    defparam i10_2_lut_rep_253.init = 16'h6666;
    LUT4 LessThan_1430_i12_3_lut_3_lut (.A(n7895[7]), .B(count_c[7]), .C(n10), 
         .Z(n12)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    defparam LessThan_1430_i12_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_4_lut (.A(\reset_count[5] ), .B(n27079), .C(\reset_count[6] ), 
         .D(\reset_count[4] ), .Z(n27080)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hfcec;
    LUT4 i1_2_lut (.A(\reset_count[8] ), .B(\reset_count[7] ), .Z(n27079)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i14133_2_lut (.A(n28[0]), .B(n8019), .Z(n42[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam i14133_2_lut.init = 16'h2222;
    LUT4 i2262_4_lut (.A(n28893), .B(n25195), .C(n30647), .D(n27223), 
         .Z(n8019)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam i2262_4_lut.init = 16'ha0a8;
    LUT4 i8_4_lut (.A(n15_adj_378), .B(\count[8] ), .C(n14), .D(\count[9] ), 
         .Z(n25195)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(\count[5] ), .B(\count[6] ), .C(count[0]), .D(\count[1] ), 
         .Z(n15_adj_378)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_3_lut (.A(count[12]), .B(count_c[7]), .C(\count[3] ), .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5_3_lut.init = 16'h8080;
    LUT4 i12_4_lut (.A(count[12]), .B(n27347), .C(n20), .D(\count[1] ), 
         .Z(n10501)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i12_4_lut.init = 16'h0010;
    LUT4 i20977_4_lut (.A(count[0]), .B(n27327), .C(n27231), .D(\count[3] ), 
         .Z(n27347)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20977_4_lut.init = 16'hfffe;
    LUT4 i20957_4_lut (.A(count[11]), .B(count_c[7]), .C(\count[5] ), 
         .D(\count[9] ), .Z(n27327)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20957_4_lut.init = 16'hfffe;
    LUT4 i20865_2_lut (.A(count_c[10]), .B(\count[6] ), .Z(n27231)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20865_2_lut.init = 16'heeee;
    CCU2D add_9_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24581), .S0(n43[11]), .S1(n43[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_13.INIT0 = 16'h5aaa;
    defparam add_9_13.INIT1 = 16'h5aaa;
    defparam add_9_13.INJECT1_0 = "NO";
    defparam add_9_13.INJECT1_1 = "NO";
    CCU2D add_9_11 (.A0(\count[9] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24580), .COUT(n24581), .S0(n43[9]), .S1(n43[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_11.INIT0 = 16'h5aaa;
    defparam add_9_11.INIT1 = 16'h5aaa;
    defparam add_9_11.INJECT1_0 = "NO";
    defparam add_9_11.INJECT1_1 = "NO";
    CCU2D add_9_9 (.A0(count_c[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count[8] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24579), .COUT(n24580), .S0(n43[7]), .S1(n43[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_9.INIT0 = 16'h5aaa;
    defparam add_9_9.INIT1 = 16'h5aaa;
    defparam add_9_9.INJECT1_0 = "NO";
    defparam add_9_9.INJECT1_1 = "NO";
    CCU2D add_9_7 (.A0(\count[5] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count[6] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24578), .COUT(n24579), .S0(n43[5]), .S1(n43[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_7.INIT0 = 16'h5aaa;
    defparam add_9_7.INIT1 = 16'h5aaa;
    defparam add_9_7.INJECT1_0 = "NO";
    defparam add_9_7.INJECT1_1 = "NO";
    CCU2D add_9_5 (.A0(\count[3] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24577), .COUT(n24578), .S0(n43[3]), .S1(n43[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_5.INIT0 = 16'h5aaa;
    defparam add_9_5.INIT1 = 16'h5aaa;
    defparam add_9_5.INJECT1_0 = "NO";
    defparam add_9_5.INJECT1_1 = "NO";
    CCU2D add_9_3 (.A0(\count[1] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count[2] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24576), .COUT(n24577), .S0(n43[1]), .S1(n43[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_3.INIT0 = 16'h5aaa;
    defparam add_9_3.INIT1 = 16'h5aaa;
    defparam add_9_3.INJECT1_0 = "NO";
    defparam add_9_3.INJECT1_1 = "NO";
    CCU2D add_9_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24576), 
          .S1(n28[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_1.INIT0 = 16'hF000;
    defparam add_9_1.INIT1 = 16'h5555;
    defparam add_9_1.INJECT1_0 = "NO";
    defparam add_9_1.INJECT1_1 = "NO";
    CCU2D add_2154_9 (.A0(latched_width[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24575), .S0(n7895[7]), .S1(n7904));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2154_9.INIT0 = 16'h5555;
    defparam add_2154_9.INIT1 = 16'h0000;
    defparam add_2154_9.INJECT1_0 = "NO";
    defparam add_2154_9.INJECT1_1 = "NO";
    CCU2D add_2154_7 (.A0(latched_width[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24574), .COUT(n24575), .S0(n7898), .S1(n7897));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2154_7.INIT0 = 16'h5555;
    defparam add_2154_7.INIT1 = 16'h5555;
    defparam add_2154_7.INJECT1_0 = "NO";
    defparam add_2154_7.INJECT1_1 = "NO";
    CCU2D add_2154_5 (.A0(latched_width[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24573), .COUT(n24574), .S0(n7900), .S1(n7895[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2154_5.INIT0 = 16'h5555;
    defparam add_2154_5.INIT1 = 16'h5555;
    defparam add_2154_5.INJECT1_0 = "NO";
    defparam add_2154_5.INJECT1_1 = "NO";
    CCU2D add_2154_3 (.A0(latched_width[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24572), .COUT(n24573), .S0(n7902), .S1(n7901));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2154_3.INIT0 = 16'h5555;
    defparam add_2154_3.INIT1 = 16'h5555;
    defparam add_2154_3.INJECT1_0 = "NO";
    defparam add_2154_3.INJECT1_1 = "NO";
    CCU2D add_2154_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(latched_width[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24572), .S1(n7903));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2154_1.INIT0 = 16'hF000;
    defparam add_2154_1.INIT1 = 16'h5555;
    defparam add_2154_1.INJECT1_0 = "NO";
    defparam add_2154_1.INJECT1_1 = "NO";
    FD1P3IX latched_width_i0_i7 (.D(\register[0] [7]), .SP(n10501), .CD(n14439), 
            .CK(debug_c_c), .Q(latched_width[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i7.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i6 (.D(\register[0] [6]), .SP(n10501), .PD(n14439), 
            .CK(debug_c_c), .Q(latched_width[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i6.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i5 (.D(\register[0] [5]), .SP(n10501), .PD(n14439), 
            .CK(debug_c_c), .Q(latched_width[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i5.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i4 (.D(\register[0] [4]), .SP(n10501), .PD(n14439), 
            .CK(debug_c_c), .Q(latched_width[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i4.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i3 (.D(\register[0] [3]), .SP(n10501), .PD(n14439), 
            .CK(debug_c_c), .Q(latched_width[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i3.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i2 (.D(\register[0] [2]), .SP(n10501), .PD(n14439), 
            .CK(debug_c_c), .Q(latched_width[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i2.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i1 (.D(\register[0] [1]), .SP(n10501), .PD(n14439), 
            .CK(debug_c_c), .Q(latched_width[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i1.GSR = "ENABLED";
    OFS1P3IX pwm_19 (.D(n25126), .SP(n28893), .SCLK(debug_c_c), .CD(GND_net), 
            .Q(motor_pwm_l_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam pwm_19.GSR = "ENABLED";
    LUT4 i9_2_lut_rep_300 (.A(n7895[4]), .B(count_c[4]), .Z(n28958)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    defparam i9_2_lut_rep_300.init = 16'h6666;
    LUT4 LessThan_1430_i8_3_lut_3_lut (.A(n7895[4]), .B(count_c[4]), .C(n6), 
         .Z(n8)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    defparam LessThan_1430_i8_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_adj_466 (.A(count_c[10]), .B(n3582), .Z(n6_adj_184)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(26[9:19])
    defparam i1_2_lut_adj_466.init = 16'heeee;
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b010000) 
//

module \ArmPeripheral(axis_haddr=8'b010000)  (GND_net, n24974, stepping, 
            n14, \register_addr[0] , n15, \register_addr[1] , Stepper_Y_M0_c_0, 
            debug_c_c, n30649, VCC_net, Stepper_Y_nFault_c, \read_size[0] , 
            n26778, n580, prev_select, n28974, databus, n3359, n7840, 
            n30651, n30648, n30650, \control_reg[7] , Stepper_Y_Dir_c, 
            n30652, Stepper_Y_M2_c_2, Stepper_Y_M1_c_1, \read_size[2] , 
            n26869, n30653, \steps_reg[5] , \steps_reg[3] , n30647, 
            Stepper_Y_En_c, Stepper_Y_Step_c, n8050, read_value, n28966, 
            n28936, \register_addr[5] , limit_c_1, n28991) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n24974;
    input stepping;
    input n14;
    input \register_addr[0] ;
    input n15;
    input \register_addr[1] ;
    output Stepper_Y_M0_c_0;
    input debug_c_c;
    input n30649;
    input VCC_net;
    input Stepper_Y_nFault_c;
    output \read_size[0] ;
    input n26778;
    input n580;
    output prev_select;
    input n28974;
    input [31:0]databus;
    input n3359;
    input n7840;
    input n30651;
    input n30648;
    input n30650;
    output \control_reg[7] ;
    output Stepper_Y_Dir_c;
    input n30652;
    output Stepper_Y_M2_c_2;
    output Stepper_Y_M1_c_1;
    output \read_size[2] ;
    input n26869;
    input n30653;
    output \steps_reg[5] ;
    output \steps_reg[3] ;
    input n30647;
    output Stepper_Y_En_c;
    output Stepper_Y_Step_c;
    input n8050;
    output [31:0]read_value;
    input n28966;
    input n28936;
    input \register_addr[5] ;
    input limit_c_1;
    input n28991;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n24389;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n225;
    
    wire n24390, n49, n62, n58, n50, step_clk, prev_step_clk, 
        n18863, n18865, n18866, n18868;
    wire [7:0]n7321;
    
    wire n5;
    wire [31:0]n5464;
    
    wire n27478;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n27479;
    wire [31:0]n3360;
    
    wire fault_latched, n12916, n41, n60, n54, n42, n20621, limit_latched, 
        n183, prev_limit_latched, n12398, n52, n38, int_step, n20627, 
        n28906, n28915, n9602;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n27400, n27401, n27403, n27404, n56, n46, n26797, n26799, 
        n26807, n26808, n26809, n26810, n26811, n26806, n26798, 
        n26812, n26813, n26800, n26805, n26819, n26801, n26814, 
        n26802, n26817, n26815, n26803, n26816, n26821, n26820, 
        n26804, n26818, n27402, n27405, n27480;
    wire [31:0]n5428;
    
    wire n24404, n24403, n24402, n24401, n24400, n24399, n24398, 
        n24397, n24396, n24395, n24394, n24393, n24392, n24391;
    
    CCU2D sub_126_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24389), .COUT(n24390), .S0(n225[1]), .S1(n225[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_3.INIT0 = 16'h5555;
    defparam sub_126_add_2_3.INIT1 = 16'h5555;
    defparam sub_126_add_2_3.INJECT1_0 = "NO";
    defparam sub_126_add_2_3.INJECT1_1 = "NO";
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n24974)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    CCU2D sub_126_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(stepping), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n24389), .S1(n225[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_1.INIT0 = 16'h0000;
    defparam sub_126_add_2_1.INIT1 = 16'h5595;
    defparam sub_126_add_2_1.INJECT1_0 = "NO";
    defparam sub_126_add_2_1.INJECT1_1 = "NO";
    PFUMX i13124 (.BLUT(n18863), .ALUT(n14), .C0(\register_addr[0] ), 
          .Z(n18865));
    PFUMX i13127 (.BLUT(n18866), .ALUT(n15), .C0(\register_addr[0] ), 
          .Z(n18868));
    PFUMX i6 (.BLUT(n7321[6]), .ALUT(n5), .C0(\register_addr[1] ), .Z(n5464[6]));
    LUT4 i17_4_lut (.A(steps_reg[0]), .B(steps_reg[9]), .C(steps_reg[28]), 
         .D(steps_reg[2]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i21108_3_lut (.A(Stepper_Y_M0_c_0), .B(stepping), .C(\register_addr[0] ), 
         .Z(n27478)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21108_3_lut.init = 16'hcaca;
    LUT4 i21109_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n27479)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21109_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i0 (.D(n3360[0]), .CK(debug_c_c), .CD(n30649), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    IFS1P3DX fault_latched_179 (.D(Stepper_Y_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_179.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n26778), .SP(n12916), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    FD1P3AX control_reg_i1 (.D(n580), .SP(n20621), .CK(debug_c_c), .Q(Stepper_Y_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_176 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_176.GSR = "ENABLED";
    FD1S3AX limit_latched_177 (.D(n183), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_177.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_178 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_178.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n580), .SP(n12398), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_175 (.D(n28974), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_175.GSR = "ENABLED";
    LUT4 i26_4_lut (.A(steps_reg[25]), .B(n52), .C(n38), .D(steps_reg[26]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 mux_1357_i30_3_lut (.A(n225[29]), .B(databus[29]), .C(n3359), 
         .Z(n3360[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i30_3_lut.init = 16'hcaca;
    FD1P3AX int_step_183 (.D(n28906), .SP(n20627), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_183.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n7840), .PD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n7840), .CD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n7840), .PD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n7840), .PD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n7840), .PD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n7840), .CD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n7840), .PD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n7840), .PD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n7840), .PD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n7840), .CD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n7840), .CD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n7840), .CD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n7840), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n28915), .CD(n9602), .CK(debug_c_c), 
            .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3IX control_reg_i7 (.D(databus[6]), .SP(n28915), .CD(n30650), 
            .CK(debug_c_c), .Q(control_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n28915), .PD(n30650), 
            .CK(debug_c_c), .Q(Stepper_Y_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n28915), .CD(n30652), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n28915), .PD(n30652), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n28915), .CD(n30652), 
            .CK(debug_c_c), .Q(Stepper_Y_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n28915), .PD(n30652), 
            .CK(debug_c_c), .Q(Stepper_Y_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n26869), .SP(n12916), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3360[31]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3360[30]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3360[29]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3360[28]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3360[27]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3360[26]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3360[25]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3360[24]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3360[23]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3360[22]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3360[21]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3360[20]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3360[19]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3360[18]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3360[17]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3360[16]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3360[15]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3360[14]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3360[13]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3360[12]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3360[11]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3360[10]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3360[9]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3360[8]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3360[7]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3360[6]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3360[5]), .CK(debug_c_c), .CD(n30653), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3360[4]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3360[3]), .CK(debug_c_c), .CD(n30653), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3360[2]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3360[1]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n12398), .CD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n12398), .CD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n12398), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_248 (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .Z(n28906)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i2_3_lut_rep_248.init = 16'h0808;
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n12398), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n12398), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n12398), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n12398), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    LUT4 i14882_4_lut_4_lut (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .D(n30647), .Z(n20627)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i14882_4_lut_4_lut.init = 16'h0038;
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n12398), .CD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n12398), .CD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n12398), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n12398), .CD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n12398), .CD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n12398), .CD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n12398), .CD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n12398), .CD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n12398), .CD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n12398), .CD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n12398), .CD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 i21030_3_lut (.A(Stepper_Y_M2_c_2), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n27400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21030_3_lut.init = 16'hcaca;
    LUT4 i21031_3_lut (.A(div_factor_reg[2]), .B(steps_reg[2]), .C(\register_addr[0] ), 
         .Z(n27401)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21031_3_lut.init = 16'hcaca;
    LUT4 i21033_3_lut (.A(Stepper_Y_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n27403)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21033_3_lut.init = 16'hcaca;
    LUT4 i21034_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n27404)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21034_3_lut.init = 16'hcaca;
    LUT4 i18_4_lut (.A(steps_reg[8]), .B(steps_reg[11]), .C(steps_reg[16]), 
         .D(steps_reg[21]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[30]), .B(steps_reg[7]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[20]), .B(n56), .C(n46), .D(steps_reg[15]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[22]), .B(steps_reg[12]), .C(steps_reg[6]), 
         .D(steps_reg[18]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[14]), .B(steps_reg[19]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i8_1_lut (.A(control_reg[6]), .Z(Stepper_Y_En_c)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(44[14:29])
    defparam i8_1_lut.init = 16'h5555;
    LUT4 i21208_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_Y_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i21208_2_lut.init = 16'h9999;
    LUT4 i24_4_lut (.A(steps_reg[13]), .B(steps_reg[17]), .C(\steps_reg[5] ), 
         .D(steps_reg[31]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut (.A(div_factor_reg[31]), .B(n26797), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n26799)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i1_2_lut (.A(\register_addr[1] ), .B(n8050), .Z(n26797)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_442 (.A(div_factor_reg[30]), .B(n26797), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n26807)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_442.init = 16'hc088;
    LUT4 i1_4_lut_adj_443 (.A(div_factor_reg[29]), .B(n26797), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n26808)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_443.init = 16'hc088;
    LUT4 i1_4_lut_adj_444 (.A(div_factor_reg[28]), .B(n26797), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n26809)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_444.init = 16'hc088;
    LUT4 i14_2_lut (.A(steps_reg[23]), .B(steps_reg[29]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[27]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[10]), .B(\steps_reg[3] ), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_445 (.A(div_factor_reg[27]), .B(n26797), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n26810)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_445.init = 16'hc088;
    LUT4 i1_4_lut_adj_446 (.A(div_factor_reg[26]), .B(n26797), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n26811)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_446.init = 16'hc088;
    LUT4 i1_4_lut_adj_447 (.A(div_factor_reg[25]), .B(n26797), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n26806)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_447.init = 16'hc088;
    LUT4 i1_4_lut_adj_448 (.A(div_factor_reg[24]), .B(n26797), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n26798)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_448.init = 16'hc088;
    LUT4 i1_4_lut_adj_449 (.A(div_factor_reg[23]), .B(n26797), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n26812)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_449.init = 16'hc088;
    LUT4 i1_4_lut_adj_450 (.A(div_factor_reg[22]), .B(n26797), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n26813)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_450.init = 16'hc088;
    LUT4 i1_4_lut_adj_451 (.A(div_factor_reg[21]), .B(n26797), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n26800)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_451.init = 16'hc088;
    LUT4 i1_4_lut_adj_452 (.A(div_factor_reg[20]), .B(n26797), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n26805)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_452.init = 16'hc088;
    LUT4 i1_4_lut_adj_453 (.A(div_factor_reg[19]), .B(n26797), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n26819)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_453.init = 16'hc088;
    LUT4 mux_1357_i1_3_lut (.A(n225[0]), .B(databus[0]), .C(n3359), .Z(n3360[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_454 (.A(div_factor_reg[18]), .B(n26797), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n26801)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_454.init = 16'hc088;
    LUT4 i1_4_lut_adj_455 (.A(div_factor_reg[17]), .B(n26797), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n26814)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_455.init = 16'hc088;
    LUT4 i1_4_lut_adj_456 (.A(div_factor_reg[16]), .B(n26797), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n26802)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_456.init = 16'hc088;
    LUT4 i1_4_lut_adj_457 (.A(div_factor_reg[15]), .B(n26797), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n26817)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_457.init = 16'hc088;
    FD1P3AX read_value__i31 (.D(n26799), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n26807), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_458 (.A(div_factor_reg[14]), .B(n26797), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n26815)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_458.init = 16'hc088;
    LUT4 i1_4_lut_adj_459 (.A(div_factor_reg[13]), .B(n26797), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n26803)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_459.init = 16'hc088;
    LUT4 i1_4_lut_adj_460 (.A(div_factor_reg[12]), .B(n26797), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n26816)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_460.init = 16'hc088;
    LUT4 i1_4_lut_adj_461 (.A(div_factor_reg[11]), .B(n26797), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n26821)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_461.init = 16'hc088;
    LUT4 i1_4_lut_adj_462 (.A(div_factor_reg[10]), .B(n26797), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n26820)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_462.init = 16'hc088;
    FD1P3AX read_value__i29 (.D(n26808), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n26809), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_463 (.A(div_factor_reg[9]), .B(n26797), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n26804)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_463.init = 16'hc088;
    LUT4 i1_4_lut_adj_464 (.A(div_factor_reg[8]), .B(n26797), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n26818)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_464.init = 16'hc088;
    FD1P3AX read_value__i27 (.D(n26810), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n26811), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n26806), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n26798), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n26812), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n26813), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n26800), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n26805), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n26819), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n26801), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n26814), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n26802), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n26817), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    LUT4 i21248_2_lut_4_lut (.A(n28966), .B(n28936), .C(\register_addr[5] ), 
         .D(n30647), .Z(n20621)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i21248_2_lut_4_lut.init = 16'hff02;
    FD1P3AX read_value__i14 (.D(n26815), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    LUT4 mux_1357_i29_3_lut (.A(n225[28]), .B(databus[28]), .C(n3359), 
         .Z(n3360[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i29_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i13 (.D(n26803), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n26816), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n26821), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n26820), .SP(n12916), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n26804), .SP(n12916), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n26818), .SP(n12916), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n5464[7]), .SP(n12916), .CD(n8050), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    LUT4 mux_1357_i28_3_lut (.A(n225[27]), .B(databus[27]), .C(n3359), 
         .Z(n3360[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i28_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i6 (.D(n5464[6]), .SP(n12916), .CD(n8050), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    LUT4 mux_1357_i27_3_lut (.A(n225[26]), .B(databus[26]), .C(n3359), 
         .Z(n3360[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i27_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i5 (.D(n18865), .SP(n12916), .CD(n8050), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    LUT4 mux_1357_i8_3_lut (.A(n225[7]), .B(databus[7]), .C(n3359), .Z(n3360[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i8_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i4 (.D(n5464[4]), .SP(n12916), .CD(n8050), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n18868), .SP(n12916), .CD(n8050), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n27402), .SP(n12916), .CD(n8050), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n27405), .SP(n12916), .CD(n8050), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 mux_1357_i26_3_lut (.A(n225[25]), .B(databus[25]), .C(n3359), 
         .Z(n3360[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i7_3_lut (.A(n225[6]), .B(databus[6]), .C(n3359), .Z(n3360[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i25_3_lut (.A(n225[24]), .B(databus[24]), .C(n3359), 
         .Z(n3360[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i24_3_lut (.A(n225[23]), .B(databus[23]), .C(n3359), 
         .Z(n3360[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i23_3_lut (.A(n225[22]), .B(databus[22]), .C(n3359), 
         .Z(n3360[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i22_3_lut (.A(n225[21]), .B(databus[21]), .C(n3359), 
         .Z(n3360[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i6_3_lut (.A(n225[5]), .B(databus[5]), .C(n3359), .Z(n3360[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i21_3_lut (.A(n225[20]), .B(databus[20]), .C(n3359), 
         .Z(n3360[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i5_3_lut (.A(n225[4]), .B(databus[4]), .C(n3359), .Z(n3360[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i5_3_lut.init = 16'hcaca;
    PFUMX i21110 (.BLUT(n27478), .ALUT(n27479), .C0(\register_addr[1] ), 
          .Z(n27480));
    LUT4 mux_1357_i4_3_lut (.A(n225[3]), .B(databus[3]), .C(n3359), .Z(n3360[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i4_3_lut.init = 16'hcaca;
    LUT4 i119_1_lut (.A(limit_c_1), .Z(n183)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i119_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_adj_465 (.A(n7840), .B(n30647), .Z(n12398)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_465.init = 16'heeee;
    LUT4 mux_1357_i3_3_lut (.A(n225[2]), .B(databus[2]), .C(n3359), .Z(n3360[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i2_3_lut (.A(n225[1]), .B(databus[1]), .C(n3359), .Z(n3360[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i20_3_lut (.A(n225[19]), .B(databus[19]), .C(n3359), 
         .Z(n3360[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i19_3_lut (.A(n225[18]), .B(databus[18]), .C(n3359), 
         .Z(n3360[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i18_3_lut (.A(n225[17]), .B(databus[17]), .C(n3359), 
         .Z(n3360[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i18_3_lut.init = 16'hcaca;
    LUT4 i14109_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n7321[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14109_2_lut.init = 16'h2222;
    LUT4 mux_1616_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n5428[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1616_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i17_3_lut (.A(n225[16]), .B(databus[16]), .C(n3359), 
         .Z(n3360[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i17_3_lut.init = 16'hcaca;
    LUT4 i14107_2_lut (.A(\control_reg[7] ), .B(\register_addr[0] ), .Z(n7321[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14107_2_lut.init = 16'h2222;
    LUT4 mux_1357_i16_3_lut (.A(n225[15]), .B(databus[15]), .C(n3359), 
         .Z(n3360[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1616_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n5428[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1616_i8_3_lut.init = 16'hcaca;
    LUT4 i13122_3_lut (.A(Stepper_Y_Dir_c), .B(div_factor_reg[5]), .C(\register_addr[1] ), 
         .Z(n18863)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13122_3_lut.init = 16'hcaca;
    LUT4 i13125_3_lut (.A(control_reg[3]), .B(div_factor_reg[3]), .C(\register_addr[1] ), 
         .Z(n18866)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13125_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i0 (.D(n27480), .SP(n12916), .CD(n8050), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i14108_2_lut (.A(control_reg[6]), .B(\register_addr[0] ), .Z(n7321[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14108_2_lut.init = 16'h2222;
    LUT4 i5_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i5_3_lut.init = 16'hcaca;
    PFUMX mux_1620_i5 (.BLUT(n7321[4]), .ALUT(n5428[4]), .C0(\register_addr[1] ), 
          .Z(n5464[4]));
    PFUMX mux_1620_i8 (.BLUT(n7321[7]), .ALUT(n5428[7]), .C0(\register_addr[1] ), 
          .Z(n5464[7]));
    LUT4 mux_1357_i15_3_lut (.A(n225[14]), .B(databus[14]), .C(n3359), 
         .Z(n3360[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i15_3_lut.init = 16'hcaca;
    CCU2D sub_126_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24404), .S0(n225[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_33.INIT0 = 16'h5555;
    defparam sub_126_add_2_33.INIT1 = 16'h0000;
    defparam sub_126_add_2_33.INJECT1_0 = "NO";
    defparam sub_126_add_2_33.INJECT1_1 = "NO";
    LUT4 mux_1357_i14_3_lut (.A(n225[13]), .B(databus[13]), .C(n3359), 
         .Z(n3360[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i13_3_lut (.A(n225[12]), .B(databus[12]), .C(n3359), 
         .Z(n3360[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i13_3_lut.init = 16'hcaca;
    LUT4 i3841_3_lut (.A(prev_limit_latched), .B(n30647), .C(limit_latched), 
         .Z(n9602)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i3841_3_lut.init = 16'hdcdc;
    CCU2D sub_126_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24403), .COUT(n24404), .S0(n225[29]), 
          .S1(n225[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_31.INIT0 = 16'h5555;
    defparam sub_126_add_2_31.INIT1 = 16'h5555;
    defparam sub_126_add_2_31.INJECT1_0 = "NO";
    defparam sub_126_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24402), .COUT(n24403), .S0(n225[27]), 
          .S1(n225[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_29.INIT0 = 16'h5555;
    defparam sub_126_add_2_29.INIT1 = 16'h5555;
    defparam sub_126_add_2_29.INJECT1_0 = "NO";
    defparam sub_126_add_2_29.INJECT1_1 = "NO";
    PFUMX i21032 (.BLUT(n27400), .ALUT(n27401), .C0(\register_addr[1] ), 
          .Z(n27402));
    PFUMX i21035 (.BLUT(n27403), .ALUT(n27404), .C0(\register_addr[1] ), 
          .Z(n27405));
    CCU2D sub_126_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24401), .COUT(n24402), .S0(n225[25]), 
          .S1(n225[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_27.INIT0 = 16'h5555;
    defparam sub_126_add_2_27.INIT1 = 16'h5555;
    defparam sub_126_add_2_27.INJECT1_0 = "NO";
    defparam sub_126_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24400), .COUT(n24401), .S0(n225[23]), 
          .S1(n225[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_25.INIT0 = 16'h5555;
    defparam sub_126_add_2_25.INIT1 = 16'h5555;
    defparam sub_126_add_2_25.INJECT1_0 = "NO";
    defparam sub_126_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24399), .COUT(n24400), .S0(n225[21]), 
          .S1(n225[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_23.INIT0 = 16'h5555;
    defparam sub_126_add_2_23.INIT1 = 16'h5555;
    defparam sub_126_add_2_23.INJECT1_0 = "NO";
    defparam sub_126_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24398), .COUT(n24399), .S0(n225[19]), 
          .S1(n225[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_21.INIT0 = 16'h5555;
    defparam sub_126_add_2_21.INIT1 = 16'h5555;
    defparam sub_126_add_2_21.INJECT1_0 = "NO";
    defparam sub_126_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24397), .COUT(n24398), .S0(n225[17]), 
          .S1(n225[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_19.INIT0 = 16'h5555;
    defparam sub_126_add_2_19.INIT1 = 16'h5555;
    defparam sub_126_add_2_19.INJECT1_0 = "NO";
    defparam sub_126_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24396), .COUT(n24397), .S0(n225[15]), 
          .S1(n225[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_17.INIT0 = 16'h5555;
    defparam sub_126_add_2_17.INIT1 = 16'h5555;
    defparam sub_126_add_2_17.INJECT1_0 = "NO";
    defparam sub_126_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24395), .COUT(n24396), .S0(n225[13]), 
          .S1(n225[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_15.INIT0 = 16'h5555;
    defparam sub_126_add_2_15.INIT1 = 16'h5555;
    defparam sub_126_add_2_15.INJECT1_0 = "NO";
    defparam sub_126_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24394), .COUT(n24395), .S0(n225[11]), 
          .S1(n225[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_13.INIT0 = 16'h5555;
    defparam sub_126_add_2_13.INIT1 = 16'h5555;
    defparam sub_126_add_2_13.INJECT1_0 = "NO";
    defparam sub_126_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24393), .COUT(n24394), .S0(n225[9]), .S1(n225[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_11.INIT0 = 16'h5555;
    defparam sub_126_add_2_11.INIT1 = 16'h5555;
    defparam sub_126_add_2_11.INJECT1_0 = "NO";
    defparam sub_126_add_2_11.INJECT1_1 = "NO";
    LUT4 mux_1357_i12_3_lut (.A(n225[11]), .B(databus[11]), .C(n3359), 
         .Z(n3360[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i11_3_lut (.A(n225[10]), .B(databus[10]), .C(n3359), 
         .Z(n3360[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i32_3_lut (.A(n225[31]), .B(databus[31]), .C(n3359), 
         .Z(n3360[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i10_3_lut (.A(n225[9]), .B(databus[9]), .C(n3359), .Z(n3360[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1357_i9_3_lut (.A(n225[8]), .B(databus[8]), .C(n3359), .Z(n3360[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i9_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_2_lut_3_lut (.A(n28974), .B(prev_select), .C(n30647), 
         .Z(n12916)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i1_2_lut_2_lut_3_lut.init = 16'h0202;
    LUT4 i21254_3_lut_rep_257_4_lut (.A(n28974), .B(prev_select), .C(\register_addr[5] ), 
         .D(n28936), .Z(n28915)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i21254_3_lut_rep_257_4_lut.init = 16'h0002;
    CCU2D sub_126_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24392), .COUT(n24393), .S0(n225[7]), .S1(n225[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_9.INIT0 = 16'h5555;
    defparam sub_126_add_2_9.INIT1 = 16'h5555;
    defparam sub_126_add_2_9.INJECT1_0 = "NO";
    defparam sub_126_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24391), .COUT(n24392), .S0(n225[5]), .S1(n225[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_7.INIT0 = 16'h5555;
    defparam sub_126_add_2_7.INIT1 = 16'h5555;
    defparam sub_126_add_2_7.INJECT1_0 = "NO";
    defparam sub_126_add_2_7.INJECT1_1 = "NO";
    LUT4 mux_1357_i31_3_lut (.A(n225[30]), .B(databus[30]), .C(n3359), 
         .Z(n3360[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1357_i31_3_lut.init = 16'hcaca;
    CCU2D sub_126_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24390), .COUT(n24391), .S0(n225[3]), .S1(n225[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_5.INIT0 = 16'h5555;
    defparam sub_126_add_2_5.INIT1 = 16'h5555;
    defparam sub_126_add_2_5.INJECT1_0 = "NO";
    defparam sub_126_add_2_5.INJECT1_1 = "NO";
    ClockDivider_U7 step_clk_gen (.step_clk(step_clk), .debug_c_c(debug_c_c), 
            .n28991(n28991), .n30647(n30647), .GND_net(GND_net), .div_factor_reg({div_factor_reg})) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U7
//

module ClockDivider_U7 (step_clk, debug_c_c, n28991, n30647, GND_net, 
            div_factor_reg) /* synthesis syn_module_defined=1 */ ;
    output step_clk;
    input debug_c_c;
    input n28991;
    input n30647;
    input GND_net;
    input [31:0]div_factor_reg;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n6913, n6948, n28889;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n6982, n14372, n24340;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    wire [31:0]n40;
    
    wire n24339, n24338, n24337, n24336, n24335, n24334, n24120, 
        n24119, n24118, n24333, n24117, n24332, n24331, n24330, 
        n24116, n24115, n24329, n24328, n24327, n24326, n24325, 
        n24114, n24113, n24112, n24111, n24110, n24109, n24108, 
        n24107, n24106, n24105, n24104, n24103, n24102, n24101, 
        n24100, n24099, n24098, n24097, n24096, n24095, n24094, 
        n24093, n24092, n24091, n24090, n24555, n24554, n24089, 
        n24088, n24087, n24553, n24552, n24551, n24550, n24086, 
        n24085, n24084, n24083, n24082, n24549, n24548, n24081, 
        n24080, n24547, n24079, n24078, n24077, n24076, n24546, 
        n24545, n24075, n24074, n24544, n24073, n24543, n24542, 
        n24541, n24540;
    
    FD1S3IX clk_o_22 (.D(n6913), .CK(debug_c_c), .CD(n28991), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    LUT4 i954_2_lut_rep_231 (.A(n6948), .B(n30647), .Z(n28889)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i954_2_lut_rep_231.init = 16'heeee;
    FD1S3IX count_2169__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i0.GSR = "ENABLED";
    LUT4 i8606_2_lut_3_lut (.A(n6948), .B(n30647), .C(n6982), .Z(n14372)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i8606_2_lut_3_lut.init = 16'he0e0;
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24340), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24339), .COUT(n24340), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24338), .COUT(n24339), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24337), .COUT(n24338), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24336), .COUT(n24337), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24335), .COUT(n24336), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24334), .COUT(n24335), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24120), .S1(n6913));
    defparam sub_1715_add_2_33.INIT0 = 16'h5555;
    defparam sub_1715_add_2_33.INIT1 = 16'h0000;
    defparam sub_1715_add_2_33.INJECT1_0 = "NO";
    defparam sub_1715_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24119), .COUT(n24120));
    defparam sub_1715_add_2_31.INIT0 = 16'h5999;
    defparam sub_1715_add_2_31.INIT1 = 16'h5999;
    defparam sub_1715_add_2_31.INJECT1_0 = "NO";
    defparam sub_1715_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24118), .COUT(n24119));
    defparam sub_1715_add_2_29.INIT0 = 16'h5999;
    defparam sub_1715_add_2_29.INIT1 = 16'h5999;
    defparam sub_1715_add_2_29.INJECT1_0 = "NO";
    defparam sub_1715_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24333), .COUT(n24334), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24117), .COUT(n24118));
    defparam sub_1715_add_2_27.INIT0 = 16'h5999;
    defparam sub_1715_add_2_27.INIT1 = 16'h5999;
    defparam sub_1715_add_2_27.INJECT1_0 = "NO";
    defparam sub_1715_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24332), .COUT(n24333), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24331), .COUT(n24332), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24330), .COUT(n24331), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24116), .COUT(n24117));
    defparam sub_1715_add_2_25.INIT0 = 16'h5999;
    defparam sub_1715_add_2_25.INIT1 = 16'h5999;
    defparam sub_1715_add_2_25.INJECT1_0 = "NO";
    defparam sub_1715_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24115), .COUT(n24116));
    defparam sub_1715_add_2_23.INIT0 = 16'h5999;
    defparam sub_1715_add_2_23.INIT1 = 16'h5999;
    defparam sub_1715_add_2_23.INJECT1_0 = "NO";
    defparam sub_1715_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24329), .COUT(n24330), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24328), .COUT(n24329), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24327), .COUT(n24328), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24326), .COUT(n24327), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24325), .COUT(n24326), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24325), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24114), .COUT(n24115));
    defparam sub_1715_add_2_21.INIT0 = 16'h5999;
    defparam sub_1715_add_2_21.INIT1 = 16'h5999;
    defparam sub_1715_add_2_21.INJECT1_0 = "NO";
    defparam sub_1715_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24113), .COUT(n24114));
    defparam sub_1715_add_2_19.INIT0 = 16'h5999;
    defparam sub_1715_add_2_19.INIT1 = 16'h5999;
    defparam sub_1715_add_2_19.INJECT1_0 = "NO";
    defparam sub_1715_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24112), .COUT(n24113));
    defparam sub_1715_add_2_17.INIT0 = 16'h5999;
    defparam sub_1715_add_2_17.INIT1 = 16'h5999;
    defparam sub_1715_add_2_17.INJECT1_0 = "NO";
    defparam sub_1715_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24111), .COUT(n24112));
    defparam sub_1715_add_2_15.INIT0 = 16'h5999;
    defparam sub_1715_add_2_15.INIT1 = 16'h5999;
    defparam sub_1715_add_2_15.INJECT1_0 = "NO";
    defparam sub_1715_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24110), .COUT(n24111));
    defparam sub_1715_add_2_13.INIT0 = 16'h5999;
    defparam sub_1715_add_2_13.INIT1 = 16'h5999;
    defparam sub_1715_add_2_13.INJECT1_0 = "NO";
    defparam sub_1715_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24109), .COUT(n24110));
    defparam sub_1715_add_2_11.INIT0 = 16'h5999;
    defparam sub_1715_add_2_11.INIT1 = 16'h5999;
    defparam sub_1715_add_2_11.INJECT1_0 = "NO";
    defparam sub_1715_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24108), .COUT(n24109));
    defparam sub_1715_add_2_9.INIT0 = 16'h5999;
    defparam sub_1715_add_2_9.INIT1 = 16'h5999;
    defparam sub_1715_add_2_9.INJECT1_0 = "NO";
    defparam sub_1715_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24107), .COUT(n24108));
    defparam sub_1715_add_2_7.INIT0 = 16'h5999;
    defparam sub_1715_add_2_7.INIT1 = 16'h5999;
    defparam sub_1715_add_2_7.INJECT1_0 = "NO";
    defparam sub_1715_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24106), .COUT(n24107));
    defparam sub_1715_add_2_5.INIT0 = 16'h5999;
    defparam sub_1715_add_2_5.INIT1 = 16'h5999;
    defparam sub_1715_add_2_5.INJECT1_0 = "NO";
    defparam sub_1715_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24105), .COUT(n24106));
    defparam sub_1715_add_2_3.INIT0 = 16'h5999;
    defparam sub_1715_add_2_3.INIT1 = 16'h5999;
    defparam sub_1715_add_2_3.INJECT1_0 = "NO";
    defparam sub_1715_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1715_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n24105));
    defparam sub_1715_add_2_1.INIT0 = 16'h0000;
    defparam sub_1715_add_2_1.INIT1 = 16'h5999;
    defparam sub_1715_add_2_1.INJECT1_0 = "NO";
    defparam sub_1715_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24104), .S1(n6948));
    defparam sub_1717_add_2_33.INIT0 = 16'h5999;
    defparam sub_1717_add_2_33.INIT1 = 16'h0000;
    defparam sub_1717_add_2_33.INJECT1_0 = "NO";
    defparam sub_1717_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24103), .COUT(n24104));
    defparam sub_1717_add_2_31.INIT0 = 16'h5999;
    defparam sub_1717_add_2_31.INIT1 = 16'h5999;
    defparam sub_1717_add_2_31.INJECT1_0 = "NO";
    defparam sub_1717_add_2_31.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    CCU2D sub_1717_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24102), .COUT(n24103));
    defparam sub_1717_add_2_29.INIT0 = 16'h5999;
    defparam sub_1717_add_2_29.INIT1 = 16'h5999;
    defparam sub_1717_add_2_29.INJECT1_0 = "NO";
    defparam sub_1717_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24101), .COUT(n24102));
    defparam sub_1717_add_2_27.INIT0 = 16'h5999;
    defparam sub_1717_add_2_27.INIT1 = 16'h5999;
    defparam sub_1717_add_2_27.INJECT1_0 = "NO";
    defparam sub_1717_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24100), .COUT(n24101));
    defparam sub_1717_add_2_25.INIT0 = 16'h5999;
    defparam sub_1717_add_2_25.INIT1 = 16'h5999;
    defparam sub_1717_add_2_25.INJECT1_0 = "NO";
    defparam sub_1717_add_2_25.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n28889), .PD(n14372), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_1717_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24099), .COUT(n24100));
    defparam sub_1717_add_2_23.INIT0 = 16'h5999;
    defparam sub_1717_add_2_23.INIT1 = 16'h5999;
    defparam sub_1717_add_2_23.INJECT1_0 = "NO";
    defparam sub_1717_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24098), .COUT(n24099));
    defparam sub_1717_add_2_21.INIT0 = 16'h5999;
    defparam sub_1717_add_2_21.INIT1 = 16'h5999;
    defparam sub_1717_add_2_21.INJECT1_0 = "NO";
    defparam sub_1717_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24097), .COUT(n24098));
    defparam sub_1717_add_2_19.INIT0 = 16'h5999;
    defparam sub_1717_add_2_19.INIT1 = 16'h5999;
    defparam sub_1717_add_2_19.INJECT1_0 = "NO";
    defparam sub_1717_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24096), .COUT(n24097));
    defparam sub_1717_add_2_17.INIT0 = 16'h5999;
    defparam sub_1717_add_2_17.INIT1 = 16'h5999;
    defparam sub_1717_add_2_17.INJECT1_0 = "NO";
    defparam sub_1717_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24095), .COUT(n24096));
    defparam sub_1717_add_2_15.INIT0 = 16'h5999;
    defparam sub_1717_add_2_15.INIT1 = 16'h5999;
    defparam sub_1717_add_2_15.INJECT1_0 = "NO";
    defparam sub_1717_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24094), .COUT(n24095));
    defparam sub_1717_add_2_13.INIT0 = 16'h5999;
    defparam sub_1717_add_2_13.INIT1 = 16'h5999;
    defparam sub_1717_add_2_13.INJECT1_0 = "NO";
    defparam sub_1717_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24093), .COUT(n24094));
    defparam sub_1717_add_2_11.INIT0 = 16'h5999;
    defparam sub_1717_add_2_11.INIT1 = 16'h5999;
    defparam sub_1717_add_2_11.INJECT1_0 = "NO";
    defparam sub_1717_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24092), .COUT(n24093));
    defparam sub_1717_add_2_9.INIT0 = 16'h5999;
    defparam sub_1717_add_2_9.INIT1 = 16'h5999;
    defparam sub_1717_add_2_9.INJECT1_0 = "NO";
    defparam sub_1717_add_2_9.INJECT1_1 = "NO";
    FD1S3IX count_2169__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i1.GSR = "ENABLED";
    CCU2D sub_1717_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24091), .COUT(n24092));
    defparam sub_1717_add_2_7.INIT0 = 16'h5999;
    defparam sub_1717_add_2_7.INIT1 = 16'h5999;
    defparam sub_1717_add_2_7.INJECT1_0 = "NO";
    defparam sub_1717_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24090), .COUT(n24091));
    defparam sub_1717_add_2_5.INIT0 = 16'h5999;
    defparam sub_1717_add_2_5.INIT1 = 16'h5999;
    defparam sub_1717_add_2_5.INJECT1_0 = "NO";
    defparam sub_1717_add_2_5.INJECT1_1 = "NO";
    FD1S3IX count_2169__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i2.GSR = "ENABLED";
    FD1S3IX count_2169__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i3.GSR = "ENABLED";
    FD1S3IX count_2169__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i4.GSR = "ENABLED";
    FD1S3IX count_2169__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i5.GSR = "ENABLED";
    FD1S3IX count_2169__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i6.GSR = "ENABLED";
    FD1S3IX count_2169__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i7.GSR = "ENABLED";
    FD1S3IX count_2169__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i8.GSR = "ENABLED";
    FD1S3IX count_2169__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i9.GSR = "ENABLED";
    FD1S3IX count_2169__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i10.GSR = "ENABLED";
    FD1S3IX count_2169__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i11.GSR = "ENABLED";
    FD1S3IX count_2169__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i12.GSR = "ENABLED";
    FD1S3IX count_2169__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i13.GSR = "ENABLED";
    FD1S3IX count_2169__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i14.GSR = "ENABLED";
    FD1S3IX count_2169__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i15.GSR = "ENABLED";
    FD1S3IX count_2169__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i16.GSR = "ENABLED";
    FD1S3IX count_2169__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i17.GSR = "ENABLED";
    FD1S3IX count_2169__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i18.GSR = "ENABLED";
    FD1S3IX count_2169__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i19.GSR = "ENABLED";
    FD1S3IX count_2169__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i20.GSR = "ENABLED";
    FD1S3IX count_2169__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i21.GSR = "ENABLED";
    FD1S3IX count_2169__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i22.GSR = "ENABLED";
    FD1S3IX count_2169__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i23.GSR = "ENABLED";
    FD1S3IX count_2169__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i24.GSR = "ENABLED";
    FD1S3IX count_2169__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i25.GSR = "ENABLED";
    FD1S3IX count_2169__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i26.GSR = "ENABLED";
    FD1S3IX count_2169__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i27.GSR = "ENABLED";
    FD1S3IX count_2169__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i28.GSR = "ENABLED";
    FD1S3IX count_2169__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i29.GSR = "ENABLED";
    FD1S3IX count_2169__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i30.GSR = "ENABLED";
    FD1S3IX count_2169__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n28889), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169__i31.GSR = "ENABLED";
    CCU2D count_2169_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24555), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_33.INIT1 = 16'h0000;
    defparam count_2169_add_4_33.INJECT1_0 = "NO";
    defparam count_2169_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24554), .COUT(n24555), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2169_add_4_31.INJECT1_0 = "NO";
    defparam count_2169_add_4_31.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24089), .COUT(n24090));
    defparam sub_1717_add_2_3.INIT0 = 16'h5999;
    defparam sub_1717_add_2_3.INIT1 = 16'h5999;
    defparam sub_1717_add_2_3.INJECT1_0 = "NO";
    defparam sub_1717_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n24089));
    defparam sub_1717_add_2_1.INIT0 = 16'h0000;
    defparam sub_1717_add_2_1.INIT1 = 16'h5999;
    defparam sub_1717_add_2_1.INJECT1_0 = "NO";
    defparam sub_1717_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24088), .S1(n6982));
    defparam sub_1718_add_2_33.INIT0 = 16'hf555;
    defparam sub_1718_add_2_33.INIT1 = 16'h0000;
    defparam sub_1718_add_2_33.INJECT1_0 = "NO";
    defparam sub_1718_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24087), .COUT(n24088));
    defparam sub_1718_add_2_31.INIT0 = 16'hf555;
    defparam sub_1718_add_2_31.INIT1 = 16'hf555;
    defparam sub_1718_add_2_31.INJECT1_0 = "NO";
    defparam sub_1718_add_2_31.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24553), .COUT(n24554), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2169_add_4_29.INJECT1_0 = "NO";
    defparam count_2169_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24552), .COUT(n24553), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2169_add_4_27.INJECT1_0 = "NO";
    defparam count_2169_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24551), .COUT(n24552), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2169_add_4_25.INJECT1_0 = "NO";
    defparam count_2169_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24550), .COUT(n24551), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2169_add_4_23.INJECT1_0 = "NO";
    defparam count_2169_add_4_23.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24086), .COUT(n24087));
    defparam sub_1718_add_2_29.INIT0 = 16'hf555;
    defparam sub_1718_add_2_29.INIT1 = 16'hf555;
    defparam sub_1718_add_2_29.INJECT1_0 = "NO";
    defparam sub_1718_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24085), .COUT(n24086));
    defparam sub_1718_add_2_27.INIT0 = 16'hf555;
    defparam sub_1718_add_2_27.INIT1 = 16'hf555;
    defparam sub_1718_add_2_27.INJECT1_0 = "NO";
    defparam sub_1718_add_2_27.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n28889), .CD(n14372), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_1718_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24084), .COUT(n24085));
    defparam sub_1718_add_2_25.INIT0 = 16'hf555;
    defparam sub_1718_add_2_25.INIT1 = 16'hf555;
    defparam sub_1718_add_2_25.INJECT1_0 = "NO";
    defparam sub_1718_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24083), .COUT(n24084));
    defparam sub_1718_add_2_23.INIT0 = 16'hf555;
    defparam sub_1718_add_2_23.INIT1 = 16'hf555;
    defparam sub_1718_add_2_23.INJECT1_0 = "NO";
    defparam sub_1718_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24082), .COUT(n24083));
    defparam sub_1718_add_2_21.INIT0 = 16'hf555;
    defparam sub_1718_add_2_21.INIT1 = 16'hf555;
    defparam sub_1718_add_2_21.INJECT1_0 = "NO";
    defparam sub_1718_add_2_21.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24549), .COUT(n24550), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2169_add_4_21.INJECT1_0 = "NO";
    defparam count_2169_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24548), .COUT(n24549), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2169_add_4_19.INJECT1_0 = "NO";
    defparam count_2169_add_4_19.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24081), .COUT(n24082));
    defparam sub_1718_add_2_19.INIT0 = 16'hf555;
    defparam sub_1718_add_2_19.INIT1 = 16'hf555;
    defparam sub_1718_add_2_19.INJECT1_0 = "NO";
    defparam sub_1718_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24080), .COUT(n24081));
    defparam sub_1718_add_2_17.INIT0 = 16'hf555;
    defparam sub_1718_add_2_17.INIT1 = 16'hf555;
    defparam sub_1718_add_2_17.INJECT1_0 = "NO";
    defparam sub_1718_add_2_17.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24547), .COUT(n24548), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2169_add_4_17.INJECT1_0 = "NO";
    defparam count_2169_add_4_17.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24079), .COUT(n24080));
    defparam sub_1718_add_2_15.INIT0 = 16'hf555;
    defparam sub_1718_add_2_15.INIT1 = 16'hf555;
    defparam sub_1718_add_2_15.INJECT1_0 = "NO";
    defparam sub_1718_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24078), .COUT(n24079));
    defparam sub_1718_add_2_13.INIT0 = 16'hf555;
    defparam sub_1718_add_2_13.INIT1 = 16'hf555;
    defparam sub_1718_add_2_13.INJECT1_0 = "NO";
    defparam sub_1718_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24077), .COUT(n24078));
    defparam sub_1718_add_2_11.INIT0 = 16'hf555;
    defparam sub_1718_add_2_11.INIT1 = 16'hf555;
    defparam sub_1718_add_2_11.INJECT1_0 = "NO";
    defparam sub_1718_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24076), .COUT(n24077));
    defparam sub_1718_add_2_9.INIT0 = 16'hf555;
    defparam sub_1718_add_2_9.INIT1 = 16'hf555;
    defparam sub_1718_add_2_9.INJECT1_0 = "NO";
    defparam sub_1718_add_2_9.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24546), .COUT(n24547), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2169_add_4_15.INJECT1_0 = "NO";
    defparam count_2169_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24545), .COUT(n24546), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2169_add_4_13.INJECT1_0 = "NO";
    defparam count_2169_add_4_13.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24075), .COUT(n24076));
    defparam sub_1718_add_2_7.INIT0 = 16'hf555;
    defparam sub_1718_add_2_7.INIT1 = 16'hf555;
    defparam sub_1718_add_2_7.INJECT1_0 = "NO";
    defparam sub_1718_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24074), .COUT(n24075));
    defparam sub_1718_add_2_5.INIT0 = 16'hf555;
    defparam sub_1718_add_2_5.INIT1 = 16'hf555;
    defparam sub_1718_add_2_5.INJECT1_0 = "NO";
    defparam sub_1718_add_2_5.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24544), .COUT(n24545), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2169_add_4_11.INJECT1_0 = "NO";
    defparam count_2169_add_4_11.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24073), .COUT(n24074));
    defparam sub_1718_add_2_3.INIT0 = 16'hf555;
    defparam sub_1718_add_2_3.INIT1 = 16'hf555;
    defparam sub_1718_add_2_3.INJECT1_0 = "NO";
    defparam sub_1718_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1718_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n24073));
    defparam sub_1718_add_2_1.INIT0 = 16'h0000;
    defparam sub_1718_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1718_add_2_1.INJECT1_0 = "NO";
    defparam sub_1718_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24543), .COUT(n24544), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2169_add_4_9.INJECT1_0 = "NO";
    defparam count_2169_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24542), .COUT(n24543), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2169_add_4_7.INJECT1_0 = "NO";
    defparam count_2169_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24541), .COUT(n24542), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2169_add_4_5.INJECT1_0 = "NO";
    defparam count_2169_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24540), .COUT(n24541), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2169_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2169_add_4_3.INJECT1_0 = "NO";
    defparam count_2169_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2169_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24540), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2169_add_4_1.INIT0 = 16'hF000;
    defparam count_2169_add_4_1.INIT1 = 16'h0555;
    defparam count_2169_add_4_1.INJECT1_0 = "NO";
    defparam count_2169_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ProtocolInterface(baud_div=12) 
//

module \ProtocolInterface(baud_div=12)  (n28973, n29056, \read_value[22] , 
            rw, n1, debug_c_c, n30644, n1318, register_addr, n29025, 
            debug_c_7, \register_addr[1] , \steps_reg[3] , n15, \register_addr[2] , 
            n28899, n28972, n29008, n7844, n1304, n1310, \register_addr[0] , 
            n12064, databus_out, \read_value[21] , n1_adj_149, n28921, 
            n12042, n8040, databus, \read_value[20] , n1_adj_150, 
            n9, \sendcount[1] , \steps_reg[5] , n14, n29052, n30647, 
            n12230, \steps_reg[7] , n13, n11636, n28928, n29011, 
            n28990, n11618, prev_select, n28966, n53, debug_c_2, 
            \steps_reg[5]_adj_151 , n14_adj_152, debug_c_3, debug_c_4, 
            debug_c_5, n28946, prev_select_adj_153, n28910, \read_value[16] , 
            n1_adj_154, \read_value[19] , n1_adj_155, \read_value[15] , 
            n1_adj_156, \read_value[12] , n1_adj_157, \read_value[13] , 
            n1_adj_158, \read_value[1] , n1_adj_159, \read_value[18] , 
            n1_adj_160, \read_value[14] , n1_adj_161, \read_value[17] , 
            n1_adj_162, n3359, n28981, \read_value[11] , n1_adj_163, 
            \read_value[10] , n1_adj_164, \read_value[9] , n1_adj_165, 
            \read_value[8] , n1_adj_166, \read_value[31] , n1_adj_167, 
            \read_value[30] , n1_adj_168, \read_value[29] , n1_adj_169, 
            \read_value[28] , n1_adj_170, \read_value[27] , n1_adj_171, 
            n22447, \read_value[26] , n1_adj_172, \read_value[25] , 
            n1_adj_173, \read_value[24] , n1_adj_174, \steps_reg[3]_adj_175 , 
            n15_adj_176, \read_value[23] , n1_adj_177, n26939, n12590, 
            n28929, \select[4] , n28927, n29021, n27014, n14379, 
            n28937, n14380, n3176, n28974, n26870, n26869, n28917, 
            n28900, n88, n26777, n26778, n28964, n28956, n28965, 
            \steps_reg[4] , n15_adj_178, n29016, n7840, n48, \steps_reg[5]_adj_179 , 
            n14_adj_180, n84, \steps_reg[3]_adj_181 , n15_adj_182, n60, 
            n11253, n11, n9_adj_183, n10, \reg_size[2] , n29018, 
            \select[1] , n12754, \select[2] , \select[7] , n28898, 
            n3446, n4, n28936, \reset_count[14] , n26915, \reset_count[13] , 
            \reset_count[12] , \reset_count[7] , \reset_count[6] , \reset_count[5] , 
            n24690, n9387, GND_net, n9388_c) /* synthesis syn_module_defined=1 */ ;
    output n28973;
    output n29056;
    input \read_value[22] ;
    output rw;
    output n1;
    input debug_c_c;
    output n30644;
    output n1318;
    output [7:0]register_addr;
    output n29025;
    output debug_c_7;
    output \register_addr[1] ;
    input \steps_reg[3] ;
    output n15;
    output \register_addr[2] ;
    input n28899;
    output n28972;
    output n29008;
    output n7844;
    output n1304;
    output n1310;
    output \register_addr[0] ;
    input n12064;
    output [31:0]databus_out;
    input \read_value[21] ;
    output n1_adj_149;
    output n28921;
    input n12042;
    output n8040;
    input [31:0]databus;
    input \read_value[20] ;
    output n1_adj_150;
    output n9;
    output \sendcount[1] ;
    input \steps_reg[5] ;
    output n14;
    output n29052;
    input n30647;
    output n12230;
    input \steps_reg[7] ;
    output n13;
    input n11636;
    output n28928;
    output n29011;
    output n28990;
    output n11618;
    input prev_select;
    output n28966;
    output n53;
    output debug_c_2;
    input \steps_reg[5]_adj_151 ;
    output n14_adj_152;
    output debug_c_3;
    output debug_c_4;
    output debug_c_5;
    output n28946;
    input prev_select_adj_153;
    output n28910;
    input \read_value[16] ;
    output n1_adj_154;
    input \read_value[19] ;
    output n1_adj_155;
    input \read_value[15] ;
    output n1_adj_156;
    input \read_value[12] ;
    output n1_adj_157;
    input \read_value[13] ;
    output n1_adj_158;
    input \read_value[1] ;
    output n1_adj_159;
    input \read_value[18] ;
    output n1_adj_160;
    input \read_value[14] ;
    output n1_adj_161;
    input \read_value[17] ;
    output n1_adj_162;
    output n3359;
    output n28981;
    input \read_value[11] ;
    output n1_adj_163;
    input \read_value[10] ;
    output n1_adj_164;
    input \read_value[9] ;
    output n1_adj_165;
    input \read_value[8] ;
    output n1_adj_166;
    input \read_value[31] ;
    output n1_adj_167;
    input \read_value[30] ;
    output n1_adj_168;
    input \read_value[29] ;
    output n1_adj_169;
    input \read_value[28] ;
    output n1_adj_170;
    input \read_value[27] ;
    output n1_adj_171;
    output n22447;
    input \read_value[26] ;
    output n1_adj_172;
    input \read_value[25] ;
    output n1_adj_173;
    input \read_value[24] ;
    output n1_adj_174;
    input \steps_reg[3]_adj_175 ;
    output n15_adj_176;
    input \read_value[23] ;
    output n1_adj_177;
    output n26939;
    input n12590;
    output n28929;
    output \select[4] ;
    output n28927;
    output n29021;
    output n27014;
    output n14379;
    output n28937;
    output n14380;
    output n3176;
    output n28974;
    output n26870;
    output n26869;
    output n28917;
    output n28900;
    output n88;
    output n26777;
    output n26778;
    output n28964;
    output n28956;
    output n28965;
    input \steps_reg[4] ;
    output n15_adj_178;
    output n29016;
    output n7840;
    output n48;
    input \steps_reg[5]_adj_179 ;
    output n14_adj_180;
    output n84;
    input \steps_reg[3]_adj_181 ;
    output n15_adj_182;
    output n60;
    input n11253;
    input n11;
    input n9_adj_183;
    input n10;
    input \reg_size[2] ;
    input n29018;
    output \select[1] ;
    input n12754;
    output \select[2] ;
    output \select[7] ;
    input n28898;
    output n3446;
    output n4;
    output n28936;
    input \reset_count[14] ;
    input n26915;
    input \reset_count[13] ;
    input \reset_count[12] ;
    input \reset_count[7] ;
    input \reset_count[6] ;
    input \reset_count[5] ;
    output n24690;
    output n9387;
    input GND_net;
    input n9388_c;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    wire [3:0]bufcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(46[12:20])
    
    wire n29023, n28997, n2535;
    wire [31:0]n1286;
    
    wire n30646, n29085, n28952, n30641, n26710, n29026, n29885, 
        n13989;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(52[12:19])
    
    wire n28951;
    wire [7:0]n2028;
    
    wire n29887;
    wire [7:0]register_addr_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    wire [7:0]\buffer[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire escape, n28989, n29027, n29009, n7, n27099;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    
    wire n28949, n28925, n20382, n27098, n11896;
    wire [7:0]\buffer[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n11974, n24897, n24894, n24898, n24893, n24903, n25979, 
        n25967, n26065, n25969, n26055, n25955, n25971, n26057;
    wire [7:0]\buffer[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n26053, n26061, n25963, n26059, n26067, n25981, n26003, 
        n27102, n27101, n10667, n9427, n24966, n10665, n9431, 
        n1398, n1397, n1391, n26864, n26688, n10741, n26123, n26195, 
        n13354;
    wire [7:0]esc_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(51[12:20])
    
    wire n28036, n2537, n26063, n5, n26758, n24890;
    wire [7:0]n9241;
    wire [7:0]n4842;
    wire [7:0]\buffer[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]\buffer[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n4_c, n29072;
    wire [7:0]\buffer[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n29071, n29046, n29075, n26334, n29074, n29007, n29078, 
        n4_adj_274, n29077, n29047, n24731, n17, n29048, n9_adj_275, 
        n29081, n29049, n8, n8671, n9_adj_276;
    wire [4:0]n19;
    
    wire n29080, n29084, n29083, n29087;
    wire [7:0]rx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(50[13:20])
    
    wire n11509, n29051, n28933, n29086, n29090, n29089, n29093, 
        n29092, n28012, n29096, n29095, n28998, n28987, n4_adj_278, 
        n26753, n26747, n26754, n26746, n26752, n14_adj_281, n26751, 
        n8_adj_282, n4_adj_283, n6, n26755, n26756, n26757, n9329, 
        n26759, n26762, n26748, n26761, n26763, n26760, n26765, 
        n26749, n26766, n26767, n29069, n26768, n26764, n26750, 
        n26770, n26745, n26744, n11_adj_285, n26771, n29068, n26772, 
        n26773, n26775, n26769, n26774, n27245, n28919, n29010, 
        n14029, n28139, busy, n5_adj_299, n24896, n5_adj_302, n24986, 
        n5_adj_304, n24891, n5_adj_312, n24973, n5_adj_314, n24889, 
        n13_adj_315, n14391, n26685, n28416, n5_adj_316, n24888, 
        n15_adj_317, n27193, n5_adj_318, n24887, n28922, n5_adj_319, 
        n24869, n5_adj_320, n24885, n11485, send, n25036, n11221, 
        n26339, n5_adj_321, n24883, n28047, n29017, n29094, n28034, 
        n28035, n5_adj_322, n24868, n29020, n28996, n4_adj_323, 
        n29097, n4_adj_324, n4_adj_325, n29070, n4_adj_326, n29073, 
        n29082, n11609, n29019, n1687, n11_adj_327, n11_adj_328, 
        n11_adj_329, n11_adj_330, n11_adj_331, n11_adj_332, n11_adj_333, 
        n11_adj_334, n11_adj_335, n11_adj_336, n13_adj_337, n11_adj_338, 
        n8_adj_339, n11_adj_340, n11_adj_341, n11_adj_342, n11_adj_343, 
        n5_adj_344, n24857, n28944, n5_adj_345, n25008, n13988, 
        n13353;
    wire [3:0]n1682;
    
    wire n28046, n29091, n25057, n29088, n29079, n26325, n26853, 
        n26350, n5_adj_346, n25010, n5_adj_347, n25004, n5_adj_348, 
        n25002, n5_adj_349, n25001, n5_adj_350, n25018, n26349, 
        n29015, n28140, n5_adj_352, n25039, n18434, n11_adj_353, 
        n5_adj_354, n24979, n5_adj_355, n24870, n5_adj_356, n24971, 
        n7978, n24965, n24963, n24967, n24964, n5_adj_357, n5_adj_358, 
        n26707, n6_adj_359, n5_adj_360, n5_adj_361, n5_adj_362, n26795, 
        n27243, n27319, n26709, n5_adj_363, n5_adj_364, n5_adj_365, 
        n5_adj_366, n1_adj_371, n6_adj_372, n26856, n26854, n6_adj_376, 
        n1407, n6_adj_377, n26452;
    
    LUT4 Select_3581_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[22] ), 
         .D(rw), .Z(n1)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3581_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2779_2_lut_rep_365 (.A(bufcount[1]), .B(bufcount[2]), .Z(n29023)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2779_2_lut_rep_365.init = 16'heeee;
    LUT4 i2416_2_lut_rep_339_3_lut (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[3]), 
         .Z(n28997)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2416_2_lut_rep_339_3_lut.init = 16'hfefe;
    FD1P3AX rw_498_rep_410 (.D(n1286[10]), .SP(n2535), .CK(debug_c_c), 
            .Q(n30644));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498_rep_410.GSR = "ENABLED";
    FD1S3IX bufcount__i3 (.D(n29085), .CK(debug_c_c), .CD(n30646), .Q(bufcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i3.GSR = "ENABLED";
    FD1S3IX bufcount__i2 (.D(n30641), .CK(debug_c_c), .CD(n28952), .Q(bufcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i2.GSR = "ENABLED";
    LUT4 n26710_bdd_4_lut_22254 (.A(n26710), .B(n29026), .C(n1318), .D(n1286[3]), 
         .Z(n29885)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C)) */ ;
    defparam n26710_bdd_4_lut_22254.init = 16'hdd0f;
    FD1S3IX bufcount__i1 (.D(n13989), .CK(debug_c_c), .CD(n28952), .Q(bufcount[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i1.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i4 (.D(n2028[4]), .SP(n28951), .CK(debug_c_c), 
            .Q(tx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n2028[3]), .SP(n28951), .CK(debug_c_c), 
            .Q(tx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    LUT4 n26710_bdd_4_lut (.A(bufcount[1]), .B(n1286[4]), .C(bufcount[0]), 
         .D(bufcount[3]), .Z(n29887)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam n26710_bdd_4_lut.init = 16'h0080;
    FD1P3AX tx_data_i0_i1 (.D(n2028[1]), .SP(n28951), .CK(debug_c_c), 
            .Q(tx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_367 (.A(register_addr[5]), .B(register_addr[4]), .Z(n29025)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_367.init = 16'heeee;
    FD1P3AX reg_addr_i0_i7 (.D(\buffer[1] [7]), .SP(n2535), .CK(debug_c_c), 
            .Q(register_addr_c[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i7.GSR = "ENABLED";
    LUT4 i850_2_lut_rep_368 (.A(escape), .B(debug_c_7), .Z(n29026)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i850_2_lut_rep_368.init = 16'hbbbb;
    LUT4 i1_2_lut (.A(\register_addr[1] ), .B(\steps_reg[3] ), .Z(n15)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_rep_331_4_lut (.A(escape), .B(debug_c_7), .C(n26710), 
         .D(n1286[4]), .Z(n28989)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i2_3_lut_rep_331_4_lut.init = 16'hffbf;
    FD1P3AX reg_addr_i0_i6 (.D(\buffer[1] [6]), .SP(n2535), .CK(debug_c_c), 
            .Q(register_addr_c[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i6.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i5 (.D(\buffer[1] [5]), .SP(n2535), .CK(debug_c_c), 
            .Q(register_addr[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i5.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i4 (.D(\buffer[1] [4]), .SP(n2535), .CK(debug_c_c), 
            .Q(register_addr[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i4.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i3 (.D(\buffer[1] [3]), .SP(n2535), .CK(debug_c_c), 
            .Q(register_addr_c[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i3.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i2 (.D(\buffer[1] [2]), .SP(n2535), .CK(debug_c_c), 
            .Q(\register_addr[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i2.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i1 (.D(\buffer[1] [1]), .SP(n2535), .CK(debug_c_c), 
            .Q(\register_addr[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i1.GSR = "ENABLED";
    LUT4 i3_4_lut (.A(register_addr[5]), .B(n28899), .C(n28972), .D(n29008), 
         .Z(n7844)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i3_4_lut.init = 16'h0800;
    LUT4 i1_3_lut_rep_369 (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .Z(n29027)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i1_3_lut_rep_369.init = 16'hecec;
    LUT4 i2_2_lut_rep_351_4_lut (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1286[4]), .Z(n29009)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+!(D))) */ ;
    defparam i2_2_lut_rep_351_4_lut.init = 16'hecff;
    LUT4 i1_2_lut_4_lut (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1286[4]), .Z(n7)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hec00;
    LUT4 i1_2_lut_3_lut (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n27099)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut.init = 16'hfbfb;
    FD1P3IX sendcount__i0 (.D(n20382), .SP(n28949), .CD(n28925), .CK(debug_c_c), 
            .Q(sendcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i0.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_287 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n27098)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_287.init = 16'hbfbf;
    FD1S3JX state_FSM_i1 (.D(n11896), .CK(debug_c_c), .PD(n28952), .Q(n1318));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i1.GSR = "ENABLED";
    FD1P3IX buffer_0___i21 (.D(n24897), .SP(n11974), .CD(n28952), .CK(debug_c_c), 
            .Q(\buffer[2] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i21.GSR = "ENABLED";
    FD1P3IX buffer_0___i20 (.D(n24894), .SP(n11974), .CD(n28952), .CK(debug_c_c), 
            .Q(\buffer[2] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i20.GSR = "ENABLED";
    FD1P3IX buffer_0___i19 (.D(n24898), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i19.GSR = "ENABLED";
    FD1P3IX buffer_0___i18 (.D(n24893), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i18.GSR = "ENABLED";
    FD1P3IX buffer_0___i17 (.D(n24903), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i17.GSR = "ENABLED";
    FD1P3IX buffer_0___i16 (.D(n25979), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i16.GSR = "ENABLED";
    FD1P3IX buffer_0___i15 (.D(n25967), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i15.GSR = "ENABLED";
    FD1P3IX buffer_0___i14 (.D(n26065), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i14.GSR = "ENABLED";
    FD1P3IX buffer_0___i13 (.D(n25969), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i13.GSR = "ENABLED";
    FD1P3IX buffer_0___i12 (.D(n26055), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i12.GSR = "ENABLED";
    FD1P3IX buffer_0___i11 (.D(n25955), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i11.GSR = "ENABLED";
    FD1P3IX buffer_0___i10 (.D(n25971), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i10.GSR = "ENABLED";
    FD1P3IX buffer_0___i9 (.D(n26057), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i9.GSR = "ENABLED";
    FD1P3IX buffer_0___i8 (.D(n26053), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i8.GSR = "ENABLED";
    FD1P3IX buffer_0___i7 (.D(n26061), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i7.GSR = "ENABLED";
    FD1P3IX buffer_0___i6 (.D(n25963), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[0] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i6.GSR = "ENABLED";
    FD1P3IX buffer_0___i5 (.D(n26059), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[0] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i5.GSR = "ENABLED";
    FD1P3IX buffer_0___i4 (.D(n26067), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i4.GSR = "ENABLED";
    FD1P3IX buffer_0___i3 (.D(n25981), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i3.GSR = "ENABLED";
    FD1P3IX buffer_0___i2 (.D(n26003), .SP(n11974), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i2.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_288 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n27102)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_288.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_289 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n27101)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_289.init = 16'hbfbf;
    FD1S3IX state_FSM_i21 (.D(n10667), .CK(debug_c_c), .CD(n30646), .Q(n1286[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i21.GSR = "ENABLED";
    FD1S3IX state_FSM_i20 (.D(n9427), .CK(debug_c_c), .CD(n30646), .Q(n1286[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i20.GSR = "ENABLED";
    FD1S3IX state_FSM_i19 (.D(n24966), .CK(debug_c_c), .CD(n30646), .Q(n1286[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i19.GSR = "ENABLED";
    FD1S3IX state_FSM_i18 (.D(n10665), .CK(debug_c_c), .CD(n28952), .Q(n1286[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i18.GSR = "ENABLED";
    FD1S3IX state_FSM_i17 (.D(n9431), .CK(debug_c_c), .CD(n28952), .Q(n1286[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i17.GSR = "ENABLED";
    FD1S3IX state_FSM_i16 (.D(n1398), .CK(debug_c_c), .CD(n28952), .Q(n1286[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i16.GSR = "ENABLED";
    FD1S3IX state_FSM_i15 (.D(n1397), .CK(debug_c_c), .CD(n28952), .Q(n1304));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i15.GSR = "ENABLED";
    FD1S3IX state_FSM_i14 (.D(n1286[12]), .CK(debug_c_c), .CD(n28952), 
            .Q(n1286[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i14.GSR = "ENABLED";
    FD1S3IX state_FSM_i13 (.D(n1286[11]), .CK(debug_c_c), .CD(n28952), 
            .Q(n1286[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i13.GSR = "ENABLED";
    FD1S3IX state_FSM_i12 (.D(n1286[10]), .CK(debug_c_c), .CD(n28952), 
            .Q(n1286[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i12.GSR = "ENABLED";
    FD1S3IX state_FSM_i11 (.D(n1391), .CK(debug_c_c), .CD(n28952), .Q(n1286[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i11.GSR = "ENABLED";
    FD1S3IX state_FSM_i10 (.D(n1310), .CK(debug_c_c), .CD(n28952), .Q(n1286[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i10.GSR = "ENABLED";
    FD1S3IX state_FSM_i9 (.D(n1286[7]), .CK(debug_c_c), .CD(n28952), .Q(n1310));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i9.GSR = "ENABLED";
    FD1S3IX state_FSM_i8 (.D(n1286[6]), .CK(debug_c_c), .CD(n28952), .Q(n1286[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i8.GSR = "ENABLED";
    FD1S3IX state_FSM_i7 (.D(n1286[5]), .CK(debug_c_c), .CD(n28952), .Q(n1286[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i7.GSR = "ENABLED";
    FD1S3IX state_FSM_i6 (.D(n26864), .CK(debug_c_c), .CD(n28952), .Q(n1286[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i6.GSR = "ENABLED";
    FD1S3IX state_FSM_i5 (.D(n26688), .CK(debug_c_c), .CD(n28952), .Q(n1286[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i5.GSR = "ENABLED";
    FD1S3IX state_FSM_i4 (.D(n10741), .CK(debug_c_c), .CD(n28952), .Q(n1286[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i4.GSR = "ENABLED";
    FD1S3IX state_FSM_i3 (.D(n26123), .CK(debug_c_c), .CD(n28952), .Q(n1286[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i3.GSR = "ENABLED";
    FD1S3IX state_FSM_i2 (.D(n26195), .CK(debug_c_c), .CD(n28952), .Q(n1286[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i2.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i0 (.D(\buffer[1] [0]), .SP(n2535), .CK(debug_c_c), 
            .Q(\register_addr[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i0.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i0 (.D(n2028[0]), .SP(n28951), .CK(debug_c_c), 
            .Q(tx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    FD1S3IX bufcount__i0 (.D(n13354), .CK(debug_c_c), .CD(n28952), .Q(bufcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i0.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i0 (.D(n28036), .SP(n12064), .CK(debug_c_c), .Q(esc_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i0.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i0 (.D(\buffer[2] [0]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i0.GSR = "ENABLED";
    LUT4 Select_3583_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[21] ), 
         .D(rw), .Z(n1_adj_149)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3583_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_3_lut_4_lut (.A(\register_addr[1] ), .B(n28921), .C(\register_addr[0] ), 
         .D(n12042), .Z(n8040)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_4_lut.init = 16'h2000;
    FD1P3IX buffer_0___i1 (.D(n26063), .SP(n11974), .CD(n28952), .CK(debug_c_c), 
            .Q(\buffer[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i1.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(databus[9]), .B(n5), .C(n1286[13]), .D(n26758), 
         .Z(n24890)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut.init = 16'hffec;
    LUT4 Select_3585_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[20] ), 
         .D(rw), .Z(n1_adj_150)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3585_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 mux_1574_i5_3_lut (.A(n9241[4]), .B(sendcount[0]), .C(n9), .Z(n4842[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1574_i5_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_4_i4_3_lut (.A(\buffer[4] [4]), .B(\buffer[5] [4]), 
         .C(sendcount[0]), .Z(n4_c)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_4_i4_3_lut.init = 16'hacac;
    LUT4 i21047_then_3_lut (.A(\buffer[0] [5]), .B(\buffer[2] [5]), .C(\sendcount[1] ), 
         .Z(n29072)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21047_then_3_lut.init = 16'hcaca;
    LUT4 i21047_else_3_lut (.A(\buffer[3] [5]), .B(\buffer[1] [5]), .C(\sendcount[1] ), 
         .Z(n29071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21047_else_3_lut.init = 16'hcaca;
    LUT4 i4_2_lut_rep_388 (.A(n1304), .B(n1286[15]), .Z(n29046)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_2_lut_rep_388.init = 16'heeee;
    LUT4 i1_4_lut_then_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(\sendcount[1] ), 
         .D(sendcount[2]), .Z(n29075)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i1_4_lut_then_4_lut.init = 16'h0001;
    LUT4 mux_1574_i3_3_lut (.A(n9241[2]), .B(sendcount[0]), .C(n9), .Z(n4842[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1574_i3_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n1304), .B(n1286[15]), .C(n1286[13]), 
         .D(n1286[12]), .Z(n26334)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_else_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(\sendcount[1] ), 
         .D(sendcount[2]), .Z(n29074)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i1_4_lut_else_4_lut.init = 16'h4001;
    LUT4 i1_2_lut_rep_349_3_lut (.A(n1304), .B(n1286[15]), .C(n1286[12]), 
         .Z(n29007)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_349_3_lut.init = 16'hfefe;
    LUT4 i21050_then_3_lut (.A(\buffer[0] [4]), .B(\buffer[2] [4]), .C(\sendcount[1] ), 
         .Z(n29078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21050_then_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_2_i4_3_lut (.A(\buffer[4] [2]), .B(\buffer[5] [2]), 
         .C(sendcount[0]), .Z(n4_adj_274)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_2_i4_3_lut.init = 16'hacac;
    LUT4 i21050_else_3_lut (.A(\buffer[3] [4]), .B(\buffer[1] [4]), .C(\sendcount[1] ), 
         .Z(n29077)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21050_else_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_389 (.A(n1286[3]), .B(n1286[19]), .Z(n29047)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_389.init = 16'heeee;
    FD1P3AX sendcount__i3 (.D(n24731), .SP(n28949), .CK(debug_c_c), .Q(sendcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i3.GSR = "ENABLED";
    FD1P3AX sendcount__i4 (.D(n17), .SP(n28949), .CK(debug_c_c), .Q(sendcount[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i4.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_390 (.A(n1286[11]), .B(n1286[9]), .Z(n29048)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_390.init = 16'heeee;
    LUT4 i3_2_lut_3_lut_4_lut (.A(n1286[11]), .B(n1286[9]), .C(n1286[19]), 
         .D(n1286[3]), .Z(n9_adj_275)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21053_then_3_lut (.A(\buffer[0] [3]), .B(\buffer[2] [3]), .C(\sendcount[1] ), 
         .Z(n29081)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21053_then_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_391 (.A(n1286[13]), .B(n1286[7]), .C(n1286[5]), 
         .Z(n29049)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_391.init = 16'hfefe;
    LUT4 i2_2_lut_4_lut (.A(n1286[13]), .B(n1286[7]), .C(n1286[5]), .D(n1286[17]), 
         .Z(n8)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_2_lut_4_lut.init = 16'hfffe;
    LUT4 i2883_2_lut_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(sendcount[2]), 
         .Z(n8671)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2883_2_lut_3_lut.init = 16'h8080;
    LUT4 i13951_3_lut_4_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(n9_adj_276), 
         .D(sendcount[2]), .Z(n19[2])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C))) */ ;
    defparam i13951_3_lut_4_lut.init = 16'h7f8f;
    LUT4 i21053_else_3_lut (.A(\buffer[3] [3]), .B(\buffer[1] [3]), .C(\sendcount[1] ), 
         .Z(n29080)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21053_else_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_290 (.A(\register_addr[1] ), .B(\steps_reg[5] ), .Z(n14)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_290.init = 16'h8888;
    LUT4 i8131_then_4_lut (.A(bufcount[3]), .B(n1318), .C(n1286[3]), .D(n1286[4]), 
         .Z(n29084)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i8131_then_4_lut.init = 16'haaa2;
    LUT4 i8131_else_4_lut (.A(bufcount[3]), .B(n1318), .C(n1286[3]), .D(n1286[4]), 
         .Z(n29083)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i8131_else_4_lut.init = 16'h0002;
    LUT4 i21056_then_3_lut (.A(\buffer[0] [2]), .B(\buffer[2] [2]), .C(\sendcount[1] ), 
         .Z(n29087)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21056_then_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_291 (.A(rx_data[1]), .B(rx_data[4]), .C(rx_data[3]), 
         .Z(n11509)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i1_2_lut_3_lut_adj_291.init = 16'h0808;
    LUT4 i1_2_lut_rep_393 (.A(register_addr[4]), .B(\register_addr[2] ), 
         .Z(n29051)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_393.init = 16'h2222;
    LUT4 i1_2_lut_rep_394 (.A(\register_addr[1] ), .B(\register_addr[0] ), 
         .Z(n29052)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_394.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_4_lut_adj_292 (.A(\register_addr[1] ), .B(\register_addr[0] ), 
         .C(n30647), .D(n28933), .Z(n12230)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_292.init = 16'hf2f0;
    LUT4 i21056_else_3_lut (.A(\buffer[3] [2]), .B(\buffer[1] [2]), .C(\sendcount[1] ), 
         .Z(n29086)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21056_else_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_rep_350_3_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), 
         .C(\register_addr[2] ), .Z(n29008)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_2_lut_rep_350_3_lut.init = 16'h0202;
    LUT4 i21059_then_3_lut (.A(\buffer[0] [1]), .B(\buffer[2] [1]), .C(\sendcount[1] ), 
         .Z(n29090)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21059_then_3_lut.init = 16'hcaca;
    LUT4 i21059_else_3_lut (.A(\buffer[3] [1]), .B(\buffer[1] [1]), .C(\sendcount[1] ), 
         .Z(n29089)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21059_else_3_lut.init = 16'hcaca;
    FD1P3IX sendcount__i2 (.D(n19[2]), .SP(n28949), .CD(n28925), .CK(debug_c_c), 
            .Q(sendcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i2.GSR = "ENABLED";
    FD1P3IX sendcount__i1 (.D(n19[1]), .SP(n28949), .CD(n28925), .CK(debug_c_c), 
            .Q(\sendcount[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i1.GSR = "ENABLED";
    LUT4 i21491_then_3_lut (.A(\buffer[0] [0]), .B(\buffer[2] [0]), .C(\sendcount[1] ), 
         .Z(n29093)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21491_then_3_lut.init = 16'hcaca;
    LUT4 i21491_else_3_lut (.A(\buffer[3] [0]), .B(\buffer[1] [0]), .C(\sendcount[1] ), 
         .Z(n29092)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21491_else_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_293 (.A(\register_addr[1] ), .B(\steps_reg[7] ), .Z(n13)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_293.init = 16'h8888;
    LUT4 rx_data_2__bdd_4_lut (.A(rx_data[2]), .B(rx_data[3]), .C(rx_data[4]), 
         .D(rx_data[1]), .Z(n28012)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D))+!B !(C+(D))))) */ ;
    defparam rx_data_2__bdd_4_lut.init = 16'h6001;
    LUT4 i21041_then_3_lut (.A(\buffer[0] [7]), .B(\buffer[2] [7]), .C(\sendcount[1] ), 
         .Z(n29096)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21041_then_3_lut.init = 16'hcaca;
    LUT4 i21041_else_3_lut (.A(\buffer[3] [7]), .B(\buffer[1] [7]), .C(\sendcount[1] ), 
         .Z(n29095)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21041_else_3_lut.init = 16'hcaca;
    LUT4 i21_2_lut_rep_270_3_lut_4_lut (.A(n11636), .B(n28998), .C(rw), 
         .D(n29056), .Z(n28928)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i21_2_lut_rep_270_3_lut_4_lut.init = 16'h0080;
    LUT4 n29885_bdd_4_lut (.A(n29885), .B(n1286[4]), .C(n29887), .D(bufcount[2]), 
         .Z(n30641)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n29885_bdd_4_lut.init = 16'heef0;
    LUT4 i1_2_lut_rep_398 (.A(register_addr_c[7]), .B(register_addr_c[3]), 
         .Z(n29056)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_398.init = 16'heeee;
    LUT4 i1_2_lut_rep_353_3_lut (.A(register_addr_c[7]), .B(register_addr_c[3]), 
         .C(register_addr_c[6]), .Z(n29011)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_353_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_314_3_lut_4_lut (.A(register_addr_c[7]), .B(register_addr_c[3]), 
         .C(register_addr[4]), .D(register_addr_c[6]), .Z(n28972)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_314_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_329_3_lut_4_lut (.A(register_addr_c[7]), .B(register_addr_c[3]), 
         .C(register_addr[5]), .D(register_addr_c[6]), .Z(n28987)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_2_lut_rep_329_3_lut_4_lut.init = 16'hffef;
    LUT4 i1_2_lut_rep_332_3_lut_4_lut (.A(register_addr_c[7]), .B(register_addr_c[3]), 
         .C(\register_addr[2] ), .D(register_addr_c[6]), .Z(n28990)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_332_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_308_4_lut (.A(n28998), .B(n29056), .C(n11618), .D(prev_select), 
         .Z(n28966)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_308_4_lut.init = 16'h0020;
    LUT4 i21_2_lut_4_lut (.A(n28998), .B(n29056), .C(n11618), .D(rw), 
         .Z(n53)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i21_2_lut_4_lut.init = 16'h2000;
    LUT4 mux_1574_i2_3_lut (.A(n9241[1]), .B(sendcount[0]), .C(n9), .Z(n4842[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1574_i2_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_1_i4_3_lut (.A(\buffer[4] [1]), .B(\buffer[5] [1]), 
         .C(sendcount[0]), .Z(n4_adj_278)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_1_i4_3_lut.init = 16'hacac;
    LUT4 i5_4_lut (.A(n9_adj_275), .B(n1286[15]), .C(n8), .D(n1286[1]), 
         .Z(debug_c_2)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i5_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_294 (.A(\register_addr[1] ), .B(\steps_reg[5]_adj_151 ), 
         .Z(n14_adj_152)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_294.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_295 (.A(n1286[3]), .B(n26710), .C(\buffer[2] [4]), 
         .Z(n26753)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_295.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_296 (.A(n1286[3]), .B(n26710), .C(\buffer[2] [3]), 
         .Z(n26747)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_296.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_297 (.A(n1286[3]), .B(n26710), .C(\buffer[2] [2]), 
         .Z(n26754)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_297.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_298 (.A(n1286[3]), .B(n26710), .C(\buffer[2] [1]), 
         .Z(n26746)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_298.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_299 (.A(n1286[3]), .B(n26710), .C(\buffer[2] [0]), 
         .Z(n26752)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_299.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_300 (.A(n1286[3]), .B(n26710), .C(n1286[13]), 
         .Z(n14_adj_281)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_300.init = 16'hf2f2;
    LUT4 i1_2_lut_3_lut_adj_301 (.A(n1286[3]), .B(n26710), .C(\buffer[2] [5]), 
         .Z(n26751)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_301.init = 16'h2020;
    LUT4 i1_4_lut (.A(n1286[2]), .B(n29046), .C(n8_adj_282), .D(n1286[18]), 
         .Z(debug_c_3)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i3_4_lut_adj_302 (.A(n29047), .B(n1286[6]), .C(n4_adj_283), .D(n1286[10]), 
         .Z(n8_adj_282)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_302.init = 16'hfffe;
    LUT4 i1_2_lut_adj_303 (.A(n1286[11]), .B(n1286[7]), .Z(n4_adj_283)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_303.init = 16'heeee;
    FD1P3AX rw_498 (.D(n1286[10]), .SP(n2535), .CK(debug_c_c), .Q(rw));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498.GSR = "ENABLED";
    LUT4 i4_4_lut (.A(n1286[6]), .B(n29007), .C(n29049), .D(n6), .Z(debug_c_4)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_304 (.A(n1286[4]), .B(n1286[20]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_304.init = 16'heeee;
    LUT4 i3_4_lut_adj_305 (.A(n1310), .B(n26334), .C(n1286[10]), .D(n29048), 
         .Z(debug_c_5)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_305.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_306 (.A(n1286[3]), .B(n26710), .C(\buffer[2] [6]), 
         .Z(n26755)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_306.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_307 (.A(n1286[3]), .B(n26710), .C(\buffer[2] [7]), 
         .Z(n26756)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_307.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_308 (.A(n1286[3]), .B(n26710), .C(\buffer[3] [0]), 
         .Z(n26757)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_308.init = 16'h2020;
    FD1S3AX escape_501 (.D(n9329), .CK(debug_c_c), .Q(escape));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam escape_501.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_309 (.A(n1286[3]), .B(n26710), .C(\buffer[3] [1]), 
         .Z(n26758)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_309.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_310 (.A(n1286[3]), .B(n26710), .C(\buffer[3] [2]), 
         .Z(n26759)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_310.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_311 (.A(n1286[3]), .B(n26710), .C(\buffer[3] [3]), 
         .Z(n26762)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_311.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_312 (.A(n1286[3]), .B(n26710), .C(\buffer[3] [4]), 
         .Z(n26748)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_312.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_313 (.A(n1286[3]), .B(n26710), .C(\buffer[3] [5]), 
         .Z(n26761)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_313.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_314 (.A(n1286[3]), .B(n26710), .C(\buffer[3] [6]), 
         .Z(n26763)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_314.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_315 (.A(n1286[3]), .B(n26710), .C(\buffer[3] [7]), 
         .Z(n26760)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_315.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_316 (.A(n1286[3]), .B(n26710), .C(\buffer[4] [0]), 
         .Z(n26765)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_316.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_317 (.A(n1286[3]), .B(n26710), .C(\buffer[4] [1]), 
         .Z(n26749)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_317.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_318 (.A(n1286[3]), .B(n26710), .C(\buffer[4] [2]), 
         .Z(n26766)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_318.init = 16'h2020;
    LUT4 i1_2_lut_rep_252_4_lut (.A(n28946), .B(rw), .C(prev_select_adj_153), 
         .D(n29052), .Z(n28910)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_252_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_adj_319 (.A(n1286[3]), .B(n26710), .C(\buffer[4] [3]), 
         .Z(n26767)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_319.init = 16'h2020;
    LUT4 i21044_then_3_lut (.A(\buffer[0] [6]), .B(\buffer[2] [6]), .C(\sendcount[1] ), 
         .Z(n29069)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21044_then_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_320 (.A(n1286[3]), .B(n26710), .C(\buffer[4] [4]), 
         .Z(n26768)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_320.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_321 (.A(n1286[3]), .B(n26710), .C(\buffer[4] [5]), 
         .Z(n26764)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_321.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_322 (.A(n1286[3]), .B(n26710), .C(\buffer[4] [6]), 
         .Z(n26750)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_322.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_323 (.A(n1286[3]), .B(n26710), .C(\buffer[4] [7]), 
         .Z(n26770)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_323.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_324 (.A(n1286[3]), .B(n26710), .C(\buffer[5] [0]), 
         .Z(n26745)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_324.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_325 (.A(n1286[3]), .B(n26710), .C(\buffer[5] [1]), 
         .Z(n26744)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_325.init = 16'h2020;
    LUT4 i1_4_lut_adj_326 (.A(n1286[4]), .B(\buffer[0] [0]), .C(n11_adj_285), 
         .D(n14_adj_281), .Z(n26063)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_326.init = 16'heca0;
    LUT4 i1_2_lut_3_lut_adj_327 (.A(n1286[3]), .B(n26710), .C(\buffer[5] [2]), 
         .Z(n26771)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_327.init = 16'h2020;
    LUT4 Select_3593_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[16] ), 
         .D(rw), .Z(n1_adj_154)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3593_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i21044_else_3_lut (.A(\buffer[3] [6]), .B(\buffer[1] [6]), .C(\sendcount[1] ), 
         .Z(n29068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21044_else_3_lut.init = 16'hcaca;
    LUT4 Select_3587_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[19] ), 
         .D(rw), .Z(n1_adj_155)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3587_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_328 (.A(n1286[3]), .B(n26710), .C(\buffer[5] [3]), 
         .Z(n26772)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_328.init = 16'h2020;
    LUT4 Select_3595_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[15] ), 
         .D(rw), .Z(n1_adj_156)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3595_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_3601_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[12] ), 
         .D(rw), .Z(n1_adj_157)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3601_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_329 (.A(n1286[3]), .B(n26710), .C(\buffer[5] [4]), 
         .Z(n26773)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_329.init = 16'h2020;
    LUT4 Select_3599_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[13] ), 
         .D(rw), .Z(n1_adj_158)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3599_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_3616_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[1] ), 
         .D(rw), .Z(n1_adj_159)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3616_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_330 (.A(n1286[3]), .B(n26710), .C(\buffer[5] [5]), 
         .Z(n26775)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_330.init = 16'h2020;
    LUT4 Select_3589_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[18] ), 
         .D(rw), .Z(n1_adj_160)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3589_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_331 (.A(n1286[3]), .B(n26710), .C(\buffer[5] [6]), 
         .Z(n26769)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_331.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_332 (.A(n1286[3]), .B(n26710), .C(\buffer[5] [7]), 
         .Z(n26774)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_332.init = 16'h2020;
    LUT4 Select_3597_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[14] ), 
         .D(rw), .Z(n1_adj_161)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3597_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_3591_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[17] ), 
         .D(rw), .Z(n1_adj_162)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3591_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i3_4_lut_adj_333 (.A(n28966), .B(n27245), .C(n28990), .D(n28919), 
         .Z(n3359)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(111[11:14])
    defparam i3_4_lut_adj_333.init = 16'h0200;
    LUT4 mux_512_i4_3_lut_4_lut (.A(n29010), .B(n1286[15]), .C(n1286[18]), 
         .D(esc_data[3]), .Z(n2028[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_512_i4_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_512_i5_3_lut_4_lut (.A(n29010), .B(n1286[15]), .C(n1286[18]), 
         .D(esc_data[4]), .Z(n2028[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_512_i5_3_lut_4_lut.init = 16'hf808;
    LUT4 i21213_2_lut_3_lut_4_lut (.A(n29010), .B(n1286[15]), .C(n1286[18]), 
         .D(n28981), .Z(n14029)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i21213_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i14856_3_lut_rep_293_4_lut (.A(n29010), .B(n1286[15]), .C(n1286[18]), 
         .D(n28981), .Z(n28951)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i14856_3_lut_rep_293_4_lut.init = 16'hf800;
    LUT4 i20879_2_lut (.A(n30644), .B(register_addr[5]), .Z(n27245)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20879_2_lut.init = 16'heeee;
    LUT4 Select_3603_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[11] ), 
         .D(rw), .Z(n1_adj_163)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3603_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_3605_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[10] ), 
         .D(rw), .Z(n1_adj_164)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3605_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 n26794_bdd_4_lut (.A(sendcount[3]), .B(sendcount[0]), .C(\sendcount[1] ), 
         .D(sendcount[2]), .Z(n28139)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam n26794_bdd_4_lut.init = 16'h4001;
    LUT4 mux_512_i2_3_lut_4_lut (.A(n29010), .B(n1286[15]), .C(n1286[18]), 
         .D(esc_data[1]), .Z(n2028[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_512_i2_3_lut_4_lut.init = 16'hf808;
    LUT4 i3670_3_lut_4_lut (.A(n29010), .B(n1286[15]), .C(busy), .D(n1286[16]), 
         .Z(n9431)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3670_3_lut_4_lut.init = 16'h8f88;
    LUT4 mux_512_i1_3_lut_4_lut (.A(n29010), .B(n1286[15]), .C(n1286[18]), 
         .D(esc_data[0]), .Z(n2028[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_512_i1_3_lut_4_lut.init = 16'hf808;
    LUT4 Select_3607_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[9] ), 
         .D(rw), .Z(n1_adj_165)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3607_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_3609_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[8] ), 
         .D(rw), .Z(n1_adj_166)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3609_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_adj_334 (.A(databus[5]), .B(n5_adj_299), .C(n1286[13]), 
         .D(n26751), .Z(n24896)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_334.init = 16'hffec;
    LUT4 select_1738_Select_21_i5_4_lut (.A(\buffer[2] [5]), .B(n1286[4]), 
         .C(rx_data[5]), .D(n27099), .Z(n5_adj_299)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_21_i5_4_lut.init = 16'h88c0;
    LUT4 Select_3563_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[31] ), 
         .D(rw), .Z(n1_adj_167)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3563_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_3565_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[30] ), 
         .D(rw), .Z(n1_adj_168)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3565_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_adj_335 (.A(databus[6]), .B(n5_adj_302), .C(n1286[13]), 
         .D(n26755), .Z(n24986)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_335.init = 16'hffec;
    LUT4 Select_3567_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[29] ), 
         .D(rw), .Z(n1_adj_169)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3567_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 select_1738_Select_22_i5_4_lut (.A(\buffer[2] [6]), .B(n1286[4]), 
         .C(rx_data[6]), .D(n27099), .Z(n5_adj_302)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_22_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_336 (.A(databus[7]), .B(n5_adj_304), .C(n1286[13]), 
         .D(n26756), .Z(n24891)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_336.init = 16'hffec;
    LUT4 select_1738_Select_23_i5_4_lut (.A(\buffer[2] [7]), .B(n1286[4]), 
         .C(rx_data[7]), .D(n27099), .Z(n5_adj_304)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_23_i5_4_lut.init = 16'h88c0;
    LUT4 Select_3569_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[28] ), 
         .D(rw), .Z(n1_adj_170)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3569_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_3571_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[27] ), 
         .D(rw), .Z(n1_adj_171)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3571_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_adj_337 (.A(\register_addr[1] ), .B(\register_addr[0] ), 
         .Z(n22447)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_337.init = 16'heeee;
    LUT4 Select_3573_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[26] ), 
         .D(rw), .Z(n1_adj_172)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3573_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_3575_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[25] ), 
         .D(rw), .Z(n1_adj_173)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3575_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 Select_3577_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[24] ), 
         .D(rw), .Z(n1_adj_174)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3577_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_adj_338 (.A(\register_addr[1] ), .B(\steps_reg[3]_adj_175 ), 
         .Z(n15_adj_176)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_338.init = 16'h8888;
    LUT4 i2_4_lut_adj_339 (.A(databus[8]), .B(n5_adj_312), .C(n1286[13]), 
         .D(n26757), .Z(n24973)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_339.init = 16'hffec;
    LUT4 select_1738_Select_24_i5_4_lut (.A(\buffer[3] [0]), .B(n1286[4]), 
         .C(rx_data[0]), .D(n27098), .Z(n5_adj_312)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_24_i5_4_lut.init = 16'h88c0;
    LUT4 Select_3579_i1_2_lut_3_lut_4_lut (.A(n28973), .B(n29056), .C(\read_value[23] ), 
         .D(rw), .Z(n1_adj_177)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam Select_3579_i1_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 select_1738_Select_25_i5_4_lut (.A(\buffer[3] [1]), .B(n1286[4]), 
         .C(rx_data[1]), .D(n27098), .Z(n5)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_25_i5_4_lut.init = 16'h88c0;
    LUT4 i1_3_lut_rep_275_4_lut (.A(n28973), .B(n29056), .C(prev_select_adj_153), 
         .D(rw), .Z(n28933)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_3_lut_rep_275_4_lut.init = 16'h0002;
    LUT4 i2_4_lut_adj_340 (.A(databus[10]), .B(n5_adj_314), .C(n1286[13]), 
         .D(n26759), .Z(n24889)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_340.init = 16'hffec;
    LUT4 select_1738_Select_26_i5_4_lut (.A(\buffer[3] [2]), .B(n1286[4]), 
         .C(rx_data[2]), .D(n27098), .Z(n5_adj_314)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_26_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_adj_341 (.A(register_addr[5]), .B(register_addr[4]), .Z(n26939)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_341.init = 16'h2222;
    LUT4 i1_4_lut_adj_342 (.A(n9), .B(n13_adj_315), .C(n28981), .D(n1304), 
         .Z(n14391)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_342.init = 16'h8000;
    LUT4 i1_4_lut_adj_343 (.A(n1286[4]), .B(debug_c_7), .C(n1286[2]), 
         .D(n26685), .Z(n26123)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_343.init = 16'heeea;
    LUT4 reduce_or_459_i1_3_lut (.A(busy), .B(n1286[13]), .C(n1286[20]), 
         .Z(n1397)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam reduce_or_459_i1_3_lut.init = 16'hdcdc;
    LUT4 i1_2_lut_rep_271_3_lut_4_lut (.A(\register_addr[2] ), .B(n29011), 
         .C(n12590), .D(n11636), .Z(n28929)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_271_3_lut_4_lut.init = 16'he0f0;
    LUT4 i1_2_lut_rep_269_3_lut_4_lut (.A(\register_addr[2] ), .B(n29011), 
         .C(n29025), .D(\select[4] ), .Z(n28927)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_269_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(\register_addr[2] ), .B(n29011), 
         .C(n29021), .D(n30647), .Z(n27014)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_4_lut_adj_344 (.A(n28921), .B(\register_addr[1] ), .C(\register_addr[0] ), 
         .D(n12042), .Z(n14379)) /* synthesis lut_function=(A (D)+!A !(B+!(C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_344.init = 16'hba00;
    LUT4 esc_data_4__bdd_4_lut_22345 (.A(esc_data[4]), .B(esc_data[2]), 
         .C(esc_data[1]), .D(esc_data[3]), .Z(n28416)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D)))+!A (B+(C+(D))))) */ ;
    defparam esc_data_4__bdd_4_lut_22345.init = 16'h2081;
    LUT4 i2_4_lut_adj_345 (.A(databus[11]), .B(n5_adj_316), .C(n1286[13]), 
         .D(n26762), .Z(n24888)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_345.init = 16'hffec;
    LUT4 i1_4_lut_adj_346 (.A(n15_adj_317), .B(n1286[3]), .C(n1318), .D(n27193), 
         .Z(n26685)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (C+!(D))+!B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_346.init = 16'h50dc;
    LUT4 i1_2_lut_rep_279_3_lut_4_lut (.A(\register_addr[2] ), .B(n29011), 
         .C(n26939), .D(\select[4] ), .Z(n28937)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_279_3_lut_4_lut.init = 16'h1000;
    LUT4 i8614_2_lut_4_lut (.A(n28921), .B(\register_addr[1] ), .C(\register_addr[0] ), 
         .D(n12042), .Z(n14380)) /* synthesis lut_function=(!(A+!(B (D)+!B !(C+!(D))))) */ ;
    defparam i8614_2_lut_4_lut.init = 16'h4500;
    LUT4 select_1738_Select_27_i5_4_lut (.A(\buffer[3] [3]), .B(n1286[4]), 
         .C(rx_data[3]), .D(n27098), .Z(n5_adj_316)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_27_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_347 (.A(databus[12]), .B(n5_adj_318), .C(n1286[13]), 
         .D(n26748), .Z(n24887)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_347.init = 16'hffec;
    LUT4 i2_3_lut_4_lut_adj_348 (.A(register_addr[4]), .B(n28922), .C(register_addr[5]), 
         .D(n28933), .Z(n3176)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(111[11:14])
    defparam i2_3_lut_4_lut_adj_348.init = 16'h8000;
    LUT4 select_1738_Select_28_i5_4_lut (.A(\buffer[3] [4]), .B(n1286[4]), 
         .C(rx_data[4]), .D(n27098), .Z(n5_adj_318)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_28_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_349 (.A(databus[13]), .B(n5_adj_319), .C(n1286[13]), 
         .D(n26761), .Z(n24869)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_349.init = 16'hffec;
    LUT4 select_1738_Select_29_i5_4_lut (.A(\buffer[3] [5]), .B(n1286[4]), 
         .C(rx_data[5]), .D(n27098), .Z(n5_adj_319)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_29_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_350 (.A(databus[14]), .B(n5_adj_320), .C(n1286[13]), 
         .D(n26763), .Z(n24885)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_350.init = 16'hffec;
    LUT4 select_1738_Select_30_i5_4_lut (.A(\buffer[3] [6]), .B(n1286[4]), 
         .C(rx_data[6]), .D(n27098), .Z(n5_adj_320)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_30_i5_4_lut.init = 16'h88c0;
    LUT4 i20829_3_lut (.A(n11485), .B(escape), .C(n15_adj_317), .Z(n27193)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i20829_3_lut.init = 16'hecec;
    FD1P3AX send_491 (.D(n11221), .SP(n25036), .CK(debug_c_c), .Q(send));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam send_491.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_351 (.A(n26339), .B(rx_data[4]), .C(rx_data[1]), 
         .D(rx_data[3]), .Z(n11485)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(139[12:17])
    defparam i2_4_lut_adj_351.init = 16'hbfff;
    LUT4 i2_3_lut (.A(n1286[19]), .B(n1286[16]), .C(n11221), .Z(n25036)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i2_3_lut.init = 16'hefef;
    LUT4 i2_4_lut_adj_352 (.A(databus[15]), .B(n5_adj_321), .C(n1286[13]), 
         .D(n26760), .Z(n24883)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_352.init = 16'hffec;
    LUT4 i21354_3_lut (.A(n28981), .B(n1286[20]), .C(n1286[17]), .Z(n11221)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i21354_3_lut.init = 16'h0202;
    LUT4 select_1738_Select_31_i5_4_lut (.A(\buffer[3] [7]), .B(n1286[4]), 
         .C(rx_data[7]), .D(n27098), .Z(n5_adj_321)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_31_i5_4_lut.init = 16'h88c0;
    LUT4 i14854_3_lut_rep_291 (.A(n1286[13]), .B(n28981), .C(n1304), .Z(n28949)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i14854_3_lut_rep_291.init = 16'hc8c8;
    LUT4 i21298_2_lut_3_lut_4_lut (.A(n1286[13]), .B(n28981), .C(n1304), 
         .D(n28047), .Z(n17)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;
    defparam i21298_2_lut_3_lut_4_lut.init = 16'hf700;
    LUT4 n28034_bdd_3_lut_4_lut (.A(sendcount[2]), .B(n29017), .C(n29094), 
         .D(n28034), .Z(n28035)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam n28034_bdd_3_lut_4_lut.init = 16'hf960;
    LUT4 i2_4_lut_adj_353 (.A(databus[16]), .B(n5_adj_322), .C(n1286[13]), 
         .D(n26765), .Z(n24868)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_353.init = 16'hffec;
    LUT4 mux_429_Mux_7_i7_4_lut_4_lut (.A(n29020), .B(n28996), .C(n4_adj_323), 
         .D(n29097), .Z(n9241[7])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_7_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_3_i4_3_lut (.A(\buffer[4] [3]), .B(\buffer[5] [3]), 
         .C(sendcount[0]), .Z(n4_adj_324)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_3_i4_3_lut.init = 16'hacac;
    LUT4 select_1738_Select_32_i5_4_lut (.A(\buffer[4] [0]), .B(n1286[4]), 
         .C(rx_data[0]), .D(n27102), .Z(n5_adj_322)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_32_i5_4_lut.init = 16'h88c0;
    LUT4 mux_429_Mux_6_i7_4_lut_4_lut (.A(n29020), .B(n28996), .C(n4_adj_325), 
         .D(n29070), .Z(n9241[6])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_6_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_5_i7_4_lut_4_lut (.A(n29020), .B(n28996), .C(n4_adj_326), 
         .D(n29073), .Z(n9241[5])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_5_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_3_i7_4_lut_4_lut (.A(n29020), .B(n28996), .C(n4_adj_324), 
         .D(n29082), .Z(n9241[3])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_3_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i21216_2_lut_rep_267_3_lut (.A(n1286[13]), .B(n28981), .C(n1304), 
         .Z(n28925)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i21216_2_lut_rep_267_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_3_lut_4_lut_adj_354 (.A(n29023), .B(bufcount[3]), .C(\buffer[0] [7]), 
         .D(n11609), .Z(n26864)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_354.init = 16'h0e00;
    LUT4 i1_2_lut_rep_288_3_lut_4_lut (.A(\register_addr[2] ), .B(n29019), 
         .C(n29056), .D(n11636), .Z(n28946)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_288_3_lut_4_lut.init = 16'h0400;
    LUT4 i3_4_lut_adj_355 (.A(rx_data[4]), .B(rx_data[3]), .C(rx_data[1]), 
         .D(n26339), .Z(n15_adj_317)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(139[12:17])
    defparam i3_4_lut_adj_355.init = 16'hfffe;
    LUT4 i498_2_lut (.A(n1286[3]), .B(n1286[4]), .Z(n1687)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i498_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_rep_316_4_lut (.A(\register_addr[2] ), .B(n29019), .C(n11618), 
         .D(n29056), .Z(n28974)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_316_4_lut.init = 16'h0040;
    LUT4 i24_3_lut_4_lut (.A(bufcount[0]), .B(n29023), .C(\buffer[0] [7]), 
         .D(rx_data[7]), .Z(n11_adj_327)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_356 (.A(bufcount[0]), .B(n29023), .C(rx_data[6]), 
         .D(\buffer[0] [6]), .Z(n11_adj_328)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_356.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_357 (.A(bufcount[0]), .B(n29023), .C(\buffer[0] [5]), 
         .D(rx_data[5]), .Z(n11_adj_329)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_357.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_358 (.A(bufcount[0]), .B(n29023), .C(\buffer[0] [4]), 
         .D(rx_data[4]), .Z(n11_adj_330)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_358.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_359 (.A(bufcount[0]), .B(n29023), .C(rx_data[3]), 
         .D(\buffer[0] [3]), .Z(n11_adj_331)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_359.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_360 (.A(bufcount[0]), .B(n29023), .C(\buffer[0] [2]), 
         .D(rx_data[2]), .Z(n11_adj_332)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_360.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_361 (.A(bufcount[0]), .B(n29023), .C(\buffer[0] [1]), 
         .D(rx_data[1]), .Z(n11_adj_333)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_361.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_362 (.A(bufcount[0]), .B(n29023), .C(rx_data[0]), 
         .D(\buffer[0] [0]), .Z(n11_adj_285)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_362.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_363 (.A(bufcount[0]), .B(n29023), .C(\buffer[1] [7]), 
         .D(rx_data[7]), .Z(n11_adj_334)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_363.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_364 (.A(bufcount[0]), .B(n29023), .C(\buffer[1] [6]), 
         .D(rx_data[6]), .Z(n11_adj_335)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_364.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_365 (.A(bufcount[0]), .B(n29023), .C(rx_data[5]), 
         .D(\buffer[1] [5]), .Z(n11_adj_336)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_365.init = 16'hfd20;
    LUT4 i2_4_lut_adj_366 (.A(n13_adj_337), .B(rx_data[5]), .C(rx_data[2]), 
         .D(rx_data[0]), .Z(n26339)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(139[12:17])
    defparam i2_4_lut_adj_366.init = 16'hfeff;
    LUT4 i24_3_lut_4_lut_adj_367 (.A(bufcount[0]), .B(n29023), .C(\buffer[1] [4]), 
         .D(rx_data[4]), .Z(n11_adj_338)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_367.init = 16'hf2d0;
    LUT4 mux_429_Mux_5_i4_3_lut (.A(\buffer[4] [5]), .B(\buffer[5] [5]), 
         .C(sendcount[0]), .Z(n4_adj_326)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_5_i4_3_lut.init = 16'hacac;
    LUT4 i1_4_lut_adj_368 (.A(n28997), .B(debug_c_7), .C(n11609), .D(n8_adj_339), 
         .Z(n26195)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_368.init = 16'hdc50;
    LUT4 i24_3_lut_4_lut_adj_369 (.A(bufcount[0]), .B(n29023), .C(rx_data[3]), 
         .D(\buffer[1] [3]), .Z(n11_adj_340)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_369.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_370 (.A(bufcount[0]), .B(n29023), .C(\buffer[1] [2]), 
         .D(rx_data[2]), .Z(n11_adj_341)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_370.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_371 (.A(bufcount[0]), .B(n29023), .C(\buffer[1] [1]), 
         .D(rx_data[1]), .Z(n11_adj_342)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_371.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_372 (.A(bufcount[0]), .B(n29023), .C(rx_data[0]), 
         .D(\buffer[1] [0]), .Z(n11_adj_343)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_372.init = 16'hfd20;
    LUT4 i2_4_lut_adj_373 (.A(databus[17]), .B(n5_adj_344), .C(n1286[13]), 
         .D(n26749), .Z(n24857)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_373.init = 16'hffec;
    LUT4 i1_2_lut_3_lut_4_lut_adj_374 (.A(\register_addr[1] ), .B(n29051), 
         .C(n29011), .D(register_addr[5]), .Z(n26870)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_374.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_375 (.A(\register_addr[1] ), .B(n29051), 
         .C(register_addr[5]), .D(n29011), .Z(n26869)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_375.init = 16'h0008;
    LUT4 select_1738_Select_33_i5_4_lut (.A(\buffer[4] [1]), .B(n1286[4]), 
         .C(rx_data[1]), .D(n27102), .Z(n5_adj_344)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_33_i5_4_lut.init = 16'h88c0;
    LUT4 i1_3_lut_rep_259_4_lut (.A(\register_addr[2] ), .B(n28944), .C(\register_addr[0] ), 
         .D(\register_addr[1] ), .Z(n28917)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_3_lut_rep_259_4_lut.init = 16'heefe;
    LUT4 i2_4_lut_adj_376 (.A(databus[18]), .B(n5_adj_345), .C(n1286[13]), 
         .D(n26766), .Z(n25008)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_376.init = 16'hffec;
    LUT4 i14122_2_lut (.A(bufcount[1]), .B(n1318), .Z(n13988)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14122_2_lut.init = 16'h2222;
    LUT4 select_1738_Select_34_i5_4_lut (.A(\buffer[4] [2]), .B(n1286[4]), 
         .C(rx_data[2]), .D(n27102), .Z(n5_adj_345)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_34_i5_4_lut.init = 16'h88c0;
    LUT4 i14092_2_lut (.A(bufcount[0]), .B(n1318), .Z(n13353)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14092_2_lut.init = 16'h2222;
    PFUMX i8223 (.BLUT(n13988), .ALUT(n1682[1]), .C0(n1687), .Z(n13989));
    LUT4 sendcount_4__bdd_3_lut_21503 (.A(sendcount[4]), .B(n28046), .C(sendcount[3]), 
         .Z(n28047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam sendcount_4__bdd_3_lut_21503.init = 16'hcaca;
    LUT4 sendcount_4__bdd_4_lut_21524 (.A(sendcount[4]), .B(sendcount[0]), 
         .C(sendcount[2]), .D(\sendcount[1] ), .Z(n28046)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;
    defparam sendcount_4__bdd_4_lut_21524.init = 16'h6aaa;
    LUT4 mux_429_Mux_6_i4_3_lut (.A(\buffer[4] [6]), .B(\buffer[5] [6]), 
         .C(sendcount[0]), .Z(n4_adj_325)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_6_i4_3_lut.init = 16'hacac;
    LUT4 mux_429_Mux_1_i7_4_lut_4_lut (.A(n29020), .B(n28996), .C(n4_adj_278), 
         .D(n29091), .Z(n9241[1])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_1_i7_4_lut_4_lut.init = 16'hdc10;
    PFUMX i7588 (.BLUT(n13353), .ALUT(n25057), .C0(n1687), .Z(n13354));
    LUT4 i20835_2_lut_rep_242_3_lut_4_lut (.A(\register_addr[2] ), .B(n28944), 
         .C(rw), .D(\register_addr[1] ), .Z(n28900)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i20835_2_lut_rep_242_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_429_Mux_2_i7_4_lut_4_lut (.A(n29020), .B(n28996), .C(n4_adj_274), 
         .D(n29088), .Z(n9241[2])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_2_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i1_2_lut_adj_377 (.A(register_addr[4]), .B(register_addr[5]), .Z(n11618)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_377.init = 16'h2222;
    LUT4 mux_429_Mux_4_i7_4_lut_4_lut (.A(n29020), .B(n28996), .C(n4_c), 
         .D(n29079), .Z(n9241[4])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_4_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i21376_2_lut_3_lut_4_lut (.A(\register_addr[2] ), .B(n28944), .C(\register_addr[0] ), 
         .D(\register_addr[1] ), .Z(n88)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i21376_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_adj_378 (.A(n1286[4]), .B(n29027), .C(bufcount[0]), 
         .D(n28989), .Z(n25057)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_adj_378.init = 16'hd222;
    LUT4 reduce_or_453_i1_3_lut_4_lut (.A(n28997), .B(n11609), .C(\buffer[0] [7]), 
         .D(n1286[9]), .Z(n1391)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(158[15] 160[18])
    defparam reduce_or_453_i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i1_3_lut (.A(n15_adj_317), .B(n1286[1]), .C(n1318), .Z(n8_adj_339)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut.init = 16'hecec;
    LUT4 i1_2_lut_3_lut_4_lut_adj_379 (.A(\register_addr[1] ), .B(n29051), 
         .C(n29011), .D(register_addr[5]), .Z(n26777)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_379.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_380 (.A(\register_addr[1] ), .B(n29051), 
         .C(register_addr[5]), .D(n29011), .Z(n26778)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_380.init = 16'h0004;
    LUT4 n28416_bdd_2_lut_rep_352 (.A(n28416), .B(n26325), .Z(n29010)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n28416_bdd_2_lut_rep_352.init = 16'h2222;
    LUT4 i1_2_lut_rep_286_3_lut_4_lut (.A(register_addr_c[6]), .B(n29056), 
         .C(register_addr[5]), .D(register_addr[4]), .Z(n28944)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_286_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_306_3_lut_4_lut (.A(register_addr_c[6]), .B(n29056), 
         .C(\select[4] ), .D(\register_addr[2] ), .Z(n28964)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_306_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_298_3_lut_4_lut (.A(register_addr_c[6]), .B(n29056), 
         .C(n11636), .D(\register_addr[2] ), .Z(n28956)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_2_lut_rep_298_3_lut_4_lut.init = 16'hffef;
    LUT4 i2_3_lut_4_lut_adj_381 (.A(\buffer[0] [1]), .B(n26853), .C(\buffer[0] [0]), 
         .D(\buffer[0] [2]), .Z(n26350)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i2_3_lut_4_lut_adj_381.init = 16'h0040;
    LUT4 i2_4_lut_adj_382 (.A(databus[19]), .B(n5_adj_346), .C(n1286[13]), 
         .D(n26767), .Z(n25010)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_382.init = 16'hffec;
    LUT4 select_1738_Select_35_i5_4_lut (.A(\buffer[4] [3]), .B(n1286[4]), 
         .C(rx_data[3]), .D(n27102), .Z(n5_adj_346)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_35_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_307_3_lut_4_lut (.A(register_addr_c[6]), .B(n29056), 
         .C(n22447), .D(\register_addr[2] ), .Z(n28965)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_307_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_383 (.A(databus[20]), .B(n5_adj_347), .C(n1286[13]), 
         .D(n26768), .Z(n25004)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_383.init = 16'hffec;
    LUT4 select_1738_Select_36_i5_4_lut (.A(\buffer[4] [4]), .B(n1286[4]), 
         .C(rx_data[4]), .D(n27102), .Z(n5_adj_347)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_36_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_384 (.A(databus[21]), .B(n5_adj_348), .C(n1286[13]), 
         .D(n26764), .Z(n25002)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_384.init = 16'hffec;
    LUT4 select_1738_Select_37_i5_4_lut (.A(\buffer[4] [5]), .B(n1286[4]), 
         .C(rx_data[5]), .D(n27102), .Z(n5_adj_348)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_37_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_385 (.A(databus[22]), .B(n5_adj_349), .C(n1286[13]), 
         .D(n26750), .Z(n25001)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_385.init = 16'hffec;
    LUT4 select_1738_Select_38_i5_4_lut (.A(\buffer[4] [6]), .B(n1286[4]), 
         .C(rx_data[6]), .D(n27102), .Z(n5_adj_349)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_38_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_386 (.A(databus[23]), .B(n5_adj_350), .C(n1286[13]), 
         .D(n26770), .Z(n25018)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_386.init = 16'hffec;
    LUT4 i1_2_lut_adj_387 (.A(\register_addr[1] ), .B(\steps_reg[4] ), .Z(n15_adj_178)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_387.init = 16'h8888;
    LUT4 i2_3_lut_4_lut_adj_388 (.A(\buffer[0] [1]), .B(n26853), .C(\buffer[0] [0]), 
         .D(\buffer[0] [2]), .Z(n26349)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_4_lut_adj_388.init = 16'h0400;
    LUT4 select_1738_Select_39_i5_4_lut (.A(\buffer[4] [7]), .B(n1286[4]), 
         .C(rx_data[7]), .D(n27102), .Z(n5_adj_350)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_39_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_357 (.A(n1304), .B(sendcount[4]), .Z(n29015)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_357.init = 16'h2222;
    LUT4 expansion5_c_bdd_2_lut_21547_3_lut (.A(n1304), .B(sendcount[4]), 
         .C(n28139), .Z(n28140)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam expansion5_c_bdd_2_lut_21547_3_lut.init = 16'h2020;
    LUT4 i2_4_lut_adj_389 (.A(databus[24]), .B(n5_adj_352), .C(n1286[13]), 
         .D(n26745), .Z(n25039)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_389.init = 16'hffec;
    LUT4 i1_2_lut_rep_358 (.A(n1286[6]), .B(n1286[11]), .Z(n29016)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_358.init = 16'heeee;
    FD1P3AX databus_out_i0_i31 (.D(\buffer[5] [7]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i31.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i30 (.D(\buffer[5] [6]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i30.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i29 (.D(\buffer[5] [5]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i29.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i28 (.D(\buffer[5] [4]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i28.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i27 (.D(\buffer[5] [3]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i27.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i26 (.D(\buffer[5] [2]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i26.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i25 (.D(\buffer[5] [1]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i25.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i24 (.D(\buffer[5] [0]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i24.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i23 (.D(\buffer[4] [7]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i23.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i22 (.D(\buffer[4] [6]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i22.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i21 (.D(\buffer[4] [5]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i21.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i20 (.D(\buffer[4] [4]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i20.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i19 (.D(\buffer[4] [3]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i19.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i18 (.D(\buffer[4] [2]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i18.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i17 (.D(\buffer[4] [1]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i17.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i16 (.D(\buffer[4] [0]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i16.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i15 (.D(\buffer[3] [7]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i15.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i14 (.D(\buffer[3] [6]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i14.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i13 (.D(\buffer[3] [5]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i13.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i12 (.D(\buffer[3] [4]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i12.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i11 (.D(\buffer[3] [3]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i11.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i10 (.D(\buffer[3] [2]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i10.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i9 (.D(\buffer[3] [1]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i9.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i8 (.D(\buffer[3] [0]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i8.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i7 (.D(\buffer[2] [7]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i7.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i6 (.D(\buffer[2] [6]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i6.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i5 (.D(\buffer[2] [5]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i5.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i4 (.D(\buffer[2] [4]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i4.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i3 (.D(\buffer[2] [3]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i3.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i2 (.D(\buffer[2] [2]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i2.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i1 (.D(\buffer[2] [1]), .SP(n2537), .CK(debug_c_c), 
            .Q(databus_out[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_390 (.A(n1286[6]), .B(n1286[11]), .C(n28981), 
         .Z(n18434)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_390.init = 16'he0e0;
    FD1P3AX esc_data_i0_i4 (.D(n4842[4]), .SP(n12064), .CK(debug_c_c), 
            .Q(esc_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i4.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i2 (.D(n4842[2]), .SP(n12064), .CK(debug_c_c), 
            .Q(esc_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i2.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i1 (.D(n4842[1]), .SP(n12064), .CK(debug_c_c), 
            .Q(esc_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i1.GSR = "ENABLED";
    LUT4 select_1738_Select_40_i5_4_lut (.A(\buffer[5] [0]), .B(n1286[4]), 
         .C(rx_data[0]), .D(n27101), .Z(n5_adj_352)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_40_i5_4_lut.init = 16'h88c0;
    LUT4 i13948_2_lut_rep_359 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n29017)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13948_2_lut_rep_359.init = 16'heeee;
    LUT4 i1_2_lut_rep_338_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(sendcount[2]), 
         .Z(n28996)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam i1_2_lut_rep_338_3_lut.init = 16'h1e1e;
    LUT4 i6_4_lut (.A(n11_adj_353), .B(prev_select), .C(n27245), .D(n29008), 
         .Z(n7840)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(111[11:14])
    defparam i6_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_rep_361 (.A(\select[4] ), .B(register_addr_c[6]), .Z(n29019)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(111[11:14])
    defparam i1_2_lut_rep_361.init = 16'h2222;
    LUT4 i1_2_lut_rep_340_3_lut (.A(\select[4] ), .B(register_addr_c[6]), 
         .C(\register_addr[2] ), .Z(n28998)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(111[11:14])
    defparam i1_2_lut_rep_340_3_lut.init = 16'h0202;
    LUT4 i2_4_lut_adj_391 (.A(databus[25]), .B(n5_adj_354), .C(n1286[13]), 
         .D(n26744), .Z(n24979)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_391.init = 16'hffec;
    LUT4 i1_2_lut_rep_315_3_lut_4_lut (.A(\select[4] ), .B(register_addr_c[6]), 
         .C(n11636), .D(\register_addr[2] ), .Z(n28973)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(111[11:14])
    defparam i1_2_lut_rep_315_3_lut_4_lut.init = 16'h0020;
    LUT4 i4_3_lut_4_lut (.A(\select[4] ), .B(register_addr_c[6]), .C(register_addr[4]), 
         .D(n29056), .Z(n11_adj_353)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(111[11:14])
    defparam i4_3_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_rep_362 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n29020)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut_rep_362.init = 16'h9999;
    LUT4 select_1738_Select_41_i5_4_lut (.A(\buffer[5] [1]), .B(n1286[4]), 
         .C(rx_data[1]), .D(n27101), .Z(n5_adj_354)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_41_i5_4_lut.init = 16'h88c0;
    LUT4 n11263_bdd_4_lut_21693_4_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(\buffer[5] [0]), .D(\buffer[4] [0]), .Z(n28034)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam n11263_bdd_4_lut_21693_4_lut.init = 16'h6420;
    LUT4 i2_4_lut_adj_392 (.A(databus[26]), .B(n5_adj_355), .C(n1286[13]), 
         .D(n26771), .Z(n24870)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_392.init = 16'hffec;
    LUT4 i13952_2_lut_2_lut_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(n9_adj_276), .Z(n19[1])) /* synthesis lut_function=(!(A (B (C))+!A !(B+!(C)))) */ ;
    defparam i13952_2_lut_2_lut_3_lut.init = 16'h6f6f;
    LUT4 select_1738_Select_42_i5_4_lut (.A(\buffer[5] [2]), .B(n1286[4]), 
         .C(rx_data[2]), .D(n27101), .Z(n5_adj_355)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_42_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_393 (.A(databus[27]), .B(n5_adj_356), .C(n1286[13]), 
         .D(n26772), .Z(n24971)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_393.init = 16'hffec;
    LUT4 i1_2_lut_rep_363 (.A(\register_addr[0] ), .B(\register_addr[1] ), 
         .Z(n29021)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_363.init = 16'h8888;
    FD1P3IX buffer_0___i22 (.D(n24896), .SP(n7978), .CD(n28952), .CK(debug_c_c), 
            .Q(\buffer[2] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i22.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_261_3_lut_3_lut_4_lut (.A(\register_addr[0] ), .B(\register_addr[1] ), 
         .C(register_addr[4]), .D(n30647), .Z(n28919)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_261_3_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_264_2_lut_3_lut (.A(\register_addr[0] ), .B(\register_addr[1] ), 
         .C(n30647), .Z(n28922)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_264_2_lut_3_lut.init = 16'h0808;
    LUT4 select_1738_Select_43_i5_4_lut (.A(\buffer[5] [3]), .B(n1286[4]), 
         .C(rx_data[3]), .D(n27101), .Z(n5_adj_356)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_43_i5_4_lut.init = 16'h88c0;
    FD1P3IX buffer_0___i23 (.D(n24986), .SP(n7978), .CD(n28952), .CK(debug_c_c), 
            .Q(\buffer[2] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i23.GSR = "ENABLED";
    FD1P3IX buffer_0___i24 (.D(n24891), .SP(n7978), .CD(n28952), .CK(debug_c_c), 
            .Q(\buffer[2] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i24.GSR = "ENABLED";
    FD1P3IX buffer_0___i25 (.D(n24973), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[3] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i25.GSR = "ENABLED";
    FD1P3IX buffer_0___i26 (.D(n24890), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[3] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i26.GSR = "ENABLED";
    FD1P3IX buffer_0___i27 (.D(n24889), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[3] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i27.GSR = "ENABLED";
    FD1P3IX buffer_0___i28 (.D(n24888), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[3] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i28.GSR = "ENABLED";
    FD1P3IX buffer_0___i29 (.D(n24887), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[3] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i29.GSR = "ENABLED";
    FD1P3IX buffer_0___i30 (.D(n24869), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[3] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i30.GSR = "ENABLED";
    FD1P3IX buffer_0___i31 (.D(n24885), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[3] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i31.GSR = "ENABLED";
    FD1P3IX buffer_0___i32 (.D(n24883), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[3] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i32.GSR = "ENABLED";
    FD1P3IX buffer_0___i33 (.D(n24868), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[4] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i33.GSR = "ENABLED";
    FD1P3IX buffer_0___i34 (.D(n24857), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[4] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i34.GSR = "ENABLED";
    FD1P3IX buffer_0___i35 (.D(n25008), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[4] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i35.GSR = "ENABLED";
    FD1P3IX buffer_0___i36 (.D(n25010), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[4] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i36.GSR = "ENABLED";
    FD1P3IX buffer_0___i37 (.D(n25004), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[4] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i37.GSR = "ENABLED";
    FD1P3IX buffer_0___i38 (.D(n25002), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[4] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i38.GSR = "ENABLED";
    FD1P3IX buffer_0___i39 (.D(n25001), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[4] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i39.GSR = "ENABLED";
    FD1P3IX buffer_0___i40 (.D(n25018), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[4] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i40.GSR = "ENABLED";
    FD1P3IX buffer_0___i41 (.D(n25039), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[5] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i41.GSR = "ENABLED";
    FD1P3IX buffer_0___i42 (.D(n24979), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[5] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i42.GSR = "ENABLED";
    FD1P3IX buffer_0___i43 (.D(n24870), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[5] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i43.GSR = "ENABLED";
    FD1P3IX buffer_0___i44 (.D(n24971), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[5] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i44.GSR = "ENABLED";
    FD1P3IX buffer_0___i45 (.D(n24965), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[5] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i45.GSR = "ENABLED";
    FD1P3IX buffer_0___i46 (.D(n24963), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[5] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i46.GSR = "ENABLED";
    FD1P3IX buffer_0___i47 (.D(n24967), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[5] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i47.GSR = "ENABLED";
    FD1P3IX buffer_0___i48 (.D(n24964), .SP(n7978), .CD(n30646), .CK(debug_c_c), 
            .Q(\buffer[5] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i48.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_394 (.A(databus[28]), .B(n5_adj_357), .C(n1286[13]), 
         .D(n26773), .Z(n24965)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_394.init = 16'hffec;
    LUT4 mux_429_Mux_7_i4_3_lut (.A(\buffer[4] [7]), .B(\buffer[5] [7]), 
         .C(sendcount[0]), .Z(n4_adj_323)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_7_i4_3_lut.init = 16'hacac;
    LUT4 select_1738_Select_44_i5_4_lut (.A(\buffer[5] [4]), .B(n1286[4]), 
         .C(rx_data[4]), .D(n27101), .Z(n5_adj_357)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_44_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_395 (.A(databus[29]), .B(n5_adj_358), .C(n1286[13]), 
         .D(n26775), .Z(n24963)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_395.init = 16'hffec;
    LUT4 select_1738_Select_45_i5_4_lut (.A(\buffer[5] [5]), .B(n1286[4]), 
         .C(rx_data[5]), .D(n27101), .Z(n5_adj_358)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_45_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_396 (.A(register_addr[4]), .B(n29011), 
         .C(\register_addr[2] ), .D(register_addr[5]), .Z(n48)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_396.init = 16'hffef;
    LUT4 i4_4_lut_adj_397 (.A(rx_data[2]), .B(n26707), .C(rx_data[5]), 
         .D(n6_adj_359), .Z(n11609)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i4_4_lut_adj_397.init = 16'h0800;
    LUT4 i2_4_lut_adj_398 (.A(escape), .B(n13_adj_337), .C(debug_c_7), 
         .D(n11509), .Z(n26707)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i2_4_lut_adj_398.init = 16'h1000;
    LUT4 i2_4_lut_adj_399 (.A(databus[4]), .B(n5_adj_360), .C(n1286[13]), 
         .D(n26753), .Z(n24897)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_399.init = 16'hffec;
    LUT4 i1_2_lut_rep_263_3_lut_4_lut (.A(register_addr[4]), .B(n29011), 
         .C(\register_addr[2] ), .D(register_addr[5]), .Z(n28921)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_rep_263_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_400 (.A(databus[30]), .B(n5_adj_361), .C(n1286[13]), 
         .D(n26769), .Z(n24967)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_400.init = 16'hffec;
    LUT4 select_1738_Select_20_i5_4_lut (.A(\buffer[2] [4]), .B(n1286[4]), 
         .C(rx_data[4]), .D(n27099), .Z(n5_adj_360)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_20_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_adj_401 (.A(n1286[3]), .B(rx_data[0]), .Z(n6_adj_359)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i1_2_lut_adj_401.init = 16'h8888;
    LUT4 select_1738_Select_46_i5_4_lut (.A(\buffer[5] [6]), .B(n1286[4]), 
         .C(rx_data[6]), .D(n27101), .Z(n5_adj_361)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_46_i5_4_lut.init = 16'h88c0;
    LUT4 i21282_2_lut_2_lut (.A(n28981), .B(n7978), .Z(n11974)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i21282_2_lut_2_lut.init = 16'hdddd;
    LUT4 i2_4_lut_adj_402 (.A(n28925), .B(sendcount[3]), .C(n9_adj_276), 
         .D(n8671), .Z(n24731)) /* synthesis lut_function=(!(A+(B ((D)+!C)+!B !(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_4_lut_adj_402.init = 16'h1040;
    LUT4 i2_4_lut_adj_403 (.A(databus[31]), .B(n5_adj_362), .C(n1286[13]), 
         .D(n26774), .Z(n24964)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_403.init = 16'hffec;
    LUT4 select_1738_Select_47_i5_4_lut (.A(\buffer[5] [7]), .B(n1286[4]), 
         .C(rx_data[7]), .D(n27101), .Z(n5_adj_362)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_47_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut_adj_404 (.A(n26795), .B(debug_c_7), .C(n1318), .D(n1286[1]), 
         .Z(n11896)) /* synthesis lut_function=(A+!(B+!(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_404.init = 16'hbbba;
    LUT4 i3_4_lut_adj_405 (.A(esc_data[6]), .B(esc_data[7]), .C(esc_data[5]), 
         .D(esc_data[0]), .Z(n26325)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i3_4_lut_adj_405.init = 16'hfeff;
    LUT4 i21346_4_lut (.A(n7), .B(n27243), .C(n29026), .D(n1286[3]), 
         .Z(n7978)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C+!(D))))) */ ;
    defparam i21346_4_lut.init = 16'h0544;
    LUT4 i20877_3_lut (.A(n1286[13]), .B(n1318), .C(n1286[4]), .Z(n27243)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i20877_3_lut.init = 16'hfefe;
    LUT4 i3_4_lut_adj_406 (.A(n27319), .B(rx_data[2]), .C(rx_data[1]), 
         .D(n26709), .Z(n26710)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i3_4_lut_adj_406.init = 16'h0100;
    LUT4 i1_2_lut_adj_407 (.A(sendcount[0]), .B(sendcount[3]), .Z(n13_adj_315)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_407.init = 16'hbbbb;
    LUT4 i2_4_lut_adj_408 (.A(rx_data[4]), .B(rx_data[3]), .C(rx_data[0]), 
         .D(rx_data[1]), .Z(n26709)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_4_lut_adj_408.init = 16'h0010;
    LUT4 i880_2_lut (.A(n1286[5]), .B(n28981), .Z(n2537)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i880_2_lut.init = 16'h8888;
    LUT4 i20949_3_lut (.A(rx_data[6]), .B(rx_data[7]), .C(rx_data[5]), 
         .Z(n27319)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i20949_3_lut.init = 16'hfefe;
    LUT4 i2_4_lut_adj_409 (.A(databus[3]), .B(n5_adj_363), .C(n1286[13]), 
         .D(n26747), .Z(n24894)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_409.init = 16'hffec;
    LUT4 equal_143_i13_2_lut (.A(rx_data[6]), .B(rx_data[7]), .Z(n13_adj_337)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(139[12:17])
    defparam equal_143_i13_2_lut.init = 16'heeee;
    LUT4 select_1738_Select_19_i5_4_lut (.A(\buffer[2] [3]), .B(n1286[4]), 
         .C(rx_data[3]), .D(n27099), .Z(n5_adj_363)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_19_i5_4_lut.init = 16'h88c0;
    LUT4 i878_3_lut (.A(n1286[5]), .B(n28981), .C(n1286[10]), .Z(n2535)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i878_3_lut.init = 16'hc8c8;
    LUT4 i2_4_lut_adj_410 (.A(databus[2]), .B(n5_adj_364), .C(n1286[13]), 
         .D(n26754), .Z(n24898)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_410.init = 16'hffec;
    LUT4 select_1738_Select_18_i5_4_lut (.A(\buffer[2] [2]), .B(n1286[4]), 
         .C(rx_data[2]), .D(n27099), .Z(n5_adj_364)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_18_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_411 (.A(databus[1]), .B(n5_adj_365), .C(n1286[13]), 
         .D(n26746), .Z(n24893)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_411.init = 16'hffec;
    LUT4 select_1738_Select_17_i5_4_lut (.A(\buffer[2] [1]), .B(n1286[4]), 
         .C(rx_data[1]), .D(n27099), .Z(n5_adj_365)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_17_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_412 (.A(databus[0]), .B(n5_adj_366), .C(n1286[13]), 
         .D(n26752), .Z(n24903)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_412.init = 16'hffec;
    LUT4 select_1738_Select_16_i5_4_lut (.A(\buffer[2] [0]), .B(n1286[4]), 
         .C(rx_data[0]), .D(n27099), .Z(n5_adj_366)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1738_Select_16_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_adj_413 (.A(\register_addr[1] ), .B(\steps_reg[5]_adj_179 ), 
         .Z(n14_adj_180)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_413.init = 16'h8888;
    LUT4 i21379_2_lut_4_lut (.A(register_addr[4]), .B(n28987), .C(\register_addr[2] ), 
         .D(\register_addr[1] ), .Z(n84)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i21379_2_lut_4_lut.init = 16'h0001;
    LUT4 i1_4_lut_adj_414 (.A(n1286[4]), .B(\buffer[1] [7]), .C(n11_adj_334), 
         .D(n14_adj_281), .Z(n25979)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_414.init = 16'heca0;
    LUT4 i1_2_lut_adj_415 (.A(\register_addr[1] ), .B(\steps_reg[3]_adj_181 ), 
         .Z(n15_adj_182)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_415.init = 16'h8888;
    LUT4 i1_2_lut_4_lut_adj_416 (.A(register_addr[4]), .B(n28987), .C(\register_addr[2] ), 
         .D(\register_addr[1] ), .Z(n60)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut_adj_416.init = 16'h0100;
    LUT4 i1_4_lut_adj_417 (.A(n1286[4]), .B(\buffer[1] [6]), .C(n11_adj_335), 
         .D(n14_adj_281), .Z(n25967)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_417.init = 16'heca0;
    LUT4 i1_4_lut_adj_418 (.A(n1286[4]), .B(\buffer[1] [5]), .C(n11_adj_336), 
         .D(n14_adj_281), .Z(n26065)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_418.init = 16'heca0;
    LUT4 i1_4_lut_adj_419 (.A(n1286[4]), .B(\buffer[1] [4]), .C(n11_adj_338), 
         .D(n14_adj_281), .Z(n25969)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_419.init = 16'heca0;
    LUT4 i1_4_lut_adj_420 (.A(n1286[4]), .B(\buffer[1] [3]), .C(n11_adj_340), 
         .D(n14_adj_281), .Z(n26055)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_420.init = 16'heca0;
    LUT4 i1_4_lut_adj_421 (.A(n1286[4]), .B(\buffer[1] [2]), .C(n11_adj_341), 
         .D(n14_adj_281), .Z(n25955)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_421.init = 16'heca0;
    LUT4 i1_4_lut_adj_422 (.A(n1286[4]), .B(\buffer[1] [1]), .C(n11_adj_342), 
         .D(n14_adj_281), .Z(n25971)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_422.init = 16'heca0;
    LUT4 i1_4_lut_adj_423 (.A(n1286[4]), .B(\buffer[1] [0]), .C(n11_adj_343), 
         .D(n14_adj_281), .Z(n26057)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_423.init = 16'heca0;
    FD1P3IX esc_data_i0_i3 (.D(n9241[3]), .SP(n12064), .CD(n14391), .CK(debug_c_c), 
            .Q(esc_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i3.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i5 (.D(n9241[5]), .SP(n12064), .CD(n14391), .CK(debug_c_c), 
            .Q(esc_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i5.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i6 (.D(n9241[6]), .SP(n12064), .CD(n14391), .CK(debug_c_c), 
            .Q(esc_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i6.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i7 (.D(n9241[7]), .SP(n12064), .CD(n14391), .CK(debug_c_c), 
            .Q(esc_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i7.GSR = "ENABLED";
    LUT4 i21225_2_lut (.A(sendcount[0]), .B(n9_adj_276), .Z(n20382)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i21225_2_lut.init = 16'h7777;
    LUT4 i1_4_lut_adj_424 (.A(sendcount[4]), .B(n1_adj_371), .C(n6_adj_372), 
         .D(n11253), .Z(n9_adj_276)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i1_4_lut_adj_424.init = 16'hfeff;
    LUT4 i1_4_lut_adj_425 (.A(n1286[4]), .B(\buffer[0] [7]), .C(n11_adj_327), 
         .D(n14_adj_281), .Z(n26053)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_425.init = 16'heca0;
    LUT4 equal_48_i1_4_lut (.A(sendcount[0]), .B(n11), .C(n9_adj_183), 
         .D(n10), .Z(n1_adj_371)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam equal_48_i1_4_lut.init = 16'h5556;
    LUT4 i2_4_lut_adj_426 (.A(\reg_size[2] ), .B(sendcount[3]), .C(sendcount[2]), 
         .D(n29018), .Z(n6_adj_372)) /* synthesis lut_function=(A (B (C+!(D))+!B ((D)+!C))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i2_4_lut_adj_426.init = 16'he7de;
    LUT4 i1_4_lut_adj_427 (.A(n1286[4]), .B(\buffer[0] [6]), .C(n11_adj_328), 
         .D(n14_adj_281), .Z(n26061)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_427.init = 16'heca0;
    LUT4 i1_4_lut_adj_428 (.A(n1286[4]), .B(\buffer[0] [5]), .C(n11_adj_329), 
         .D(n14_adj_281), .Z(n25963)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_428.init = 16'heca0;
    LUT4 i2830_2_lut_3_lut_4_lut_4_lut (.A(bufcount[1]), .B(n28989), .C(n29009), 
         .D(bufcount[0]), .Z(n1682[1])) /* synthesis lut_function=(A (B (C+!(D)))+!A !((C+!(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i2830_2_lut_3_lut_4_lut_4_lut.init = 16'h8488;
    FD1P3AX select__i1 (.D(n26350), .SP(n12754), .CK(debug_c_c), .Q(\select[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i1.GSR = "ENABLED";
    FD1P3AX select__i2 (.D(n26856), .SP(n12754), .CK(debug_c_c), .Q(\select[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i2.GSR = "ENABLED";
    FD1P3AX select__i4 (.D(n26349), .SP(n12754), .CK(debug_c_c), .Q(\select[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i4.GSR = "ENABLED";
    FD1P3AX select__i7 (.D(n26854), .SP(n12754), .CK(debug_c_c), .Q(\select[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i7.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_429 (.A(n1286[4]), .B(\buffer[0] [4]), .C(n11_adj_330), 
         .D(n14_adj_281), .Z(n26059)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_429.init = 16'heca0;
    LUT4 i1_4_lut_adj_430 (.A(n1286[4]), .B(\buffer[0] [3]), .C(n11_adj_331), 
         .D(n14_adj_281), .Z(n26067)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_430.init = 16'heca0;
    FD1P3IX tx_data_i0_i2 (.D(esc_data[2]), .SP(n28951), .CD(n14029), 
            .CK(debug_c_c), .Q(tx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_431 (.A(n1286[4]), .B(\buffer[0] [2]), .C(n11_adj_332), 
         .D(n14_adj_281), .Z(n25981)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_431.init = 16'heca0;
    LUT4 i1_4_lut_adj_432 (.A(n1286[4]), .B(\buffer[0] [1]), .C(n11_adj_333), 
         .D(n14_adj_281), .Z(n26003)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_432.init = 16'heca0;
    FD1P3IX tx_data_i0_i5 (.D(esc_data[5]), .SP(n28951), .CD(n14029), 
            .CK(debug_c_c), .Q(tx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i6 (.D(esc_data[6]), .SP(n28951), .CD(n14029), 
            .CK(debug_c_c), .Q(tx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i7 (.D(esc_data[7]), .SP(n28951), .CD(n14029), 
            .CK(debug_c_c), .Q(tx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    PFUMX i21493 (.BLUT(n28035), .ALUT(n13_adj_315), .C0(n9), .Z(n28036));
    LUT4 i3_4_lut_adj_433 (.A(register_addr[5]), .B(register_addr[4]), .C(n28898), 
         .D(n27014), .Z(n3446)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i3_4_lut_adj_433.init = 16'h1000;
    LUT4 i3_4_lut_adj_434 (.A(sendcount[3]), .B(n29017), .C(sendcount[2]), 
         .D(n29015), .Z(n26795)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_434.init = 16'h0200;
    LUT4 i1_2_lut_adj_435 (.A(sendcount[0]), .B(sendcount[3]), .Z(n4)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_435.init = 16'h4444;
    LUT4 i4903_3_lut (.A(busy), .B(n1286[20]), .C(n1286[19]), .Z(n10667)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4903_3_lut.init = 16'ha8a8;
    LUT4 i2_3_lut_rep_278_4_lut (.A(n22447), .B(n28990), .C(rw), .D(register_addr[4]), 
         .Z(n28936)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_278_4_lut.init = 16'hfeff;
    LUT4 i1_4_lut_adj_436 (.A(\buffer[0] [3]), .B(n18434), .C(n6_adj_376), 
         .D(\buffer[0] [4]), .Z(n26853)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_436.init = 16'h0004;
    LUT4 i2_2_lut (.A(\buffer[0] [5]), .B(\buffer[0] [6]), .Z(n6_adj_376)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3666_3_lut (.A(n1286[19]), .B(n1286[18]), .C(busy), .Z(n9427)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3666_3_lut.init = 16'hcece;
    LUT4 i3_4_lut_adj_437 (.A(\buffer[0] [2]), .B(\buffer[0] [1]), .C(\buffer[0] [0]), 
         .D(n26853), .Z(n26856)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i3_4_lut_adj_437.init = 16'h0400;
    LUT4 i2_4_lut_adj_438 (.A(n26853), .B(\buffer[0] [0]), .C(\buffer[0] [2]), 
         .D(\buffer[0] [1]), .Z(n26854)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_4_lut_adj_438.init = 16'h8000;
    LUT4 i2_4_lut_adj_439 (.A(n29010), .B(n28140), .C(n1286[15]), .D(n1407), 
         .Z(n24966)) /* synthesis lut_function=(A (B+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_439.init = 16'hffdc;
    LUT4 i470_2_lut (.A(busy), .B(n1286[17]), .Z(n1407)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i470_2_lut.init = 16'h4444;
    LUT4 i7874_4_lut (.A(escape), .B(n11485), .C(n6_adj_377), .D(n1286[3]), 
         .Z(n9329)) /* synthesis lut_function=(!(A (C (D))+!A (B+!(C (D))))) */ ;
    defparam i7874_4_lut.init = 16'h1aaa;
    LUT4 i2_2_lut_adj_440 (.A(debug_c_7), .B(n28981), .Z(n6_adj_377)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_adj_440.init = 16'h8888;
    LUT4 i4902_3_lut (.A(busy), .B(n1286[17]), .C(n1286[16]), .Z(n10665)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4902_3_lut.init = 16'ha8a8;
    LUT4 i21295_3_lut (.A(debug_c_7), .B(n26452), .C(n1286[3]), .Z(n26688)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i21295_3_lut.init = 16'h2020;
    PFUMX i21821 (.BLUT(n29095), .ALUT(n29096), .C0(sendcount[0]), .Z(n29097));
    PFUMX i21819 (.BLUT(n29092), .ALUT(n29093), .C0(sendcount[0]), .Z(n29094));
    PFUMX i21817 (.BLUT(n29089), .ALUT(n29090), .C0(sendcount[0]), .Z(n29091));
    PFUMX i21815 (.BLUT(n29086), .ALUT(n29087), .C0(sendcount[0]), .Z(n29088));
    PFUMX i21813 (.BLUT(n29083), .ALUT(n29084), .C0(n28989), .Z(n29085));
    PFUMX i21811 (.BLUT(n29080), .ALUT(n29081), .C0(sendcount[0]), .Z(n29082));
    LUT4 i3_4_lut_adj_441 (.A(n27319), .B(n28012), .C(rx_data[0]), .D(escape), 
         .Z(n26452)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_441.init = 16'h0040;
    PFUMX i21809 (.BLUT(n29077), .ALUT(n29078), .C0(sendcount[0]), .Z(n29079));
    PFUMX i21807 (.BLUT(n29074), .ALUT(n29075), .C0(sendcount[3]), .Z(n9));
    PFUMX i21805 (.BLUT(n29071), .ALUT(n29072), .C0(sendcount[0]), .Z(n29073));
    PFUMX i21803 (.BLUT(n29068), .ALUT(n29069), .C0(sendcount[0]), .Z(n29070));
    LUT4 i461_2_lut (.A(n9), .B(n1304), .Z(n1398)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i461_2_lut.init = 16'h4444;
    \UARTTransmitter(baud_div=12)  uart_output (.\reset_count[14] (\reset_count[14] ), 
            .n26915(n26915), .\reset_count[13] (\reset_count[13] ), .\reset_count[12] (\reset_count[12] ), 
            .n30646(n30646), .n28952(n28952), .tx_data({tx_data}), .send(send), 
            .n28981(n28981), .busy(busy), .\reset_count[7] (\reset_count[7] ), 
            .\reset_count[6] (\reset_count[6] ), .\reset_count[5] (\reset_count[5] ), 
            .n24690(n24690), .n9387(n9387), .debug_c_c(debug_c_c), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(65[30] 70[52])
    \UARTReceiver(baud_div=12)  uart_input (.debug_c_7(debug_c_7), .n1315(n1286[3]), 
            .n1316(n1286[2]), .n10741(n10741), .n9388_c(n9388_c), .debug_c_c(debug_c_c), 
            .n28981(n28981), .rx_data({rx_data}), .n28952(n28952), .n30646(n30646), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(60[27] 64[39])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=12) 
//

module \UARTTransmitter(baud_div=12)  (\reset_count[14] , n26915, \reset_count[13] , 
            \reset_count[12] , n30646, n28952, tx_data, send, n28981, 
            busy, \reset_count[7] , \reset_count[6] , \reset_count[5] , 
            n24690, n9387, debug_c_c, GND_net) /* synthesis syn_module_defined=1 */ ;
    input \reset_count[14] ;
    input n26915;
    input \reset_count[13] ;
    input \reset_count[12] ;
    output n30646;
    output n28952;
    input [7:0]tx_data;
    input send;
    output n28981;
    output busy;
    input \reset_count[7] ;
    input \reset_count[6] ;
    input \reset_count[5] ;
    output n24690;
    output n9387;
    input debug_c_c;
    input GND_net;
    
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n7, n10;
    wire [3:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n104, n28001;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n7976, n28758, n28759, n12170, n25845, n17, n28000, n2529, 
        n28968, n26993, n27406, n27407, n26992, n27003, n19847, 
        n17_adj_271, n13577, n2, n27408, n27999;
    
    PFUMX Mux_22_i15 (.BLUT(n7), .ALUT(n10), .C0(state[3]), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;
    LUT4 i14853_1_lut_rep_412 (.A(\reset_count[14] ), .B(n26915), .C(\reset_count[13] ), 
         .D(\reset_count[12] ), .Z(n30646)) /* synthesis lut_function=(!(A+(B (C)+!B (C (D))))) */ ;
    defparam i14853_1_lut_rep_412.init = 16'h0515;
    FD1S3IX state__i0 (.D(n28001), .CK(bclk), .CD(n28952), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n7976), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    LUT4 state_2__bdd_4_lut_22270 (.A(state[0]), .B(state[3]), .C(state[1]), 
         .D(send), .Z(n28758)) /* synthesis lut_function=(A (B (C))+!A !(B+(C+!(D)))) */ ;
    defparam state_2__bdd_4_lut_22270.init = 16'h8180;
    LUT4 n28758_bdd_2_lut (.A(n28758), .B(state[2]), .Z(n28759)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n28758_bdd_2_lut.init = 16'h2222;
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n7976), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n7976), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n7976), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n7976), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n7976), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n7976), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n7976), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX state__i3 (.D(n25845), .SP(n12170), .CK(bclk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    LUT4 i27_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), .D(state[3]), 
         .Z(n17)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B !(C+(D))))) */ ;
    defparam i27_4_lut_4_lut.init = 16'h15fe;
    LUT4 state_1__bdd_4_lut (.A(state[1]), .B(state[3]), .C(state[0]), 
         .D(send), .Z(n28000)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(B (C)+!B (C+!(D)))) */ ;
    defparam state_1__bdd_4_lut.init = 16'h8f0e;
    LUT4 i1_2_lut (.A(state[0]), .B(state[1]), .Z(n2529)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_3_lut (.A(state[1]), .B(n28968), .C(state[0]), .Z(n26993)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4848;
    LUT4 i21036_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n27406)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21036_3_lut.init = 16'hcaca;
    LUT4 i21037_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n27407)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21037_3_lut.init = 16'hcaca;
    FD1P3AX state__i1 (.D(n26993), .SP(n12170), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    FD1P3AX state__i2 (.D(n26992), .SP(n12170), .CK(bclk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(n27003), .B(state[2]), .C(n19847), .D(n28981), 
         .Z(n7976)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i2_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_adj_286 (.A(send), .B(state[3]), .Z(n27003)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_286.init = 16'h2222;
    LUT4 i14117_2_lut (.A(state[1]), .B(state[0]), .Z(n19847)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14117_2_lut.init = 16'heeee;
    LUT4 i21363_3_lut (.A(n28981), .B(n17_adj_271), .C(state[2]), .Z(n12170)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i21363_3_lut.init = 16'hf7f7;
    LUT4 i1_4_lut (.A(n28981), .B(state[3]), .C(state[2]), .D(n2529), 
         .Z(n25845)) /* synthesis lut_function=(!((B (C)+!B !(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i1_4_lut.init = 16'h2808;
    LUT4 i3_1_lut (.A(state[3]), .Z(n13577)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i3_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_rep_323 (.A(\reset_count[14] ), .B(n26915), .C(\reset_count[13] ), 
         .D(\reset_count[12] ), .Z(n28981)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_rep_323.init = 16'hfaea;
    FD1P3IX busy_34 (.D(n13577), .SP(n28759), .CD(n30646), .CK(bclk), 
            .Q(busy));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam busy_34.GSR = "ENABLED";
    LUT4 i14853_1_lut_rep_294_4_lut (.A(\reset_count[14] ), .B(n26915), 
         .C(\reset_count[13] ), .D(\reset_count[12] ), .Z(n28952)) /* synthesis lut_function=(!(A+(B (C)+!B (C (D))))) */ ;
    defparam i14853_1_lut_rep_294_4_lut.init = 16'h0515;
    LUT4 i2_3_lut (.A(\reset_count[7] ), .B(\reset_count[6] ), .C(\reset_count[5] ), 
         .Z(n24690)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 Mux_22_i7_4_lut (.A(n2), .B(n27408), .C(state[2]), .D(state[1]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i14374_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i14374_4_lut.init = 16'hfcee;
    LUT4 state_1__bdd_2_lut (.A(state[3]), .B(state[0]), .Z(n27999)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_1__bdd_2_lut.init = 16'h1111;
    LUT4 i24_4_lut_4_lut (.A(state[3]), .B(state[0]), .C(state[1]), .D(send), 
         .Z(n17_adj_271)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;
    defparam i24_4_lut_4_lut.init = 16'h8001;
    FD1P3JX tx_35 (.D(n104), .SP(n17), .PD(n28952), .CK(bclk), .Q(n9387)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    LUT4 i1_3_lut_rep_310 (.A(n28981), .B(state[2]), .C(state[3]), .Z(n28968)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i1_3_lut_rep_310.init = 16'h2a2a;
    LUT4 i1_3_lut_4_lut (.A(n28981), .B(state[2]), .C(state[3]), .D(n2529), 
         .Z(n26992)) /* synthesis lut_function=(!((B (C+(D))+!B !(D))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h2208;
    PFUMX i21038 (.BLUT(n27406), .ALUT(n27407), .C0(state[1]), .Z(n27408));
    PFUMX i21471 (.BLUT(n28000), .ALUT(n27999), .C0(state[2]), .Z(n28001));
    \ClockDividerP(factor=12)  baud_gen (.bclk(bclk), .debug_c_c(debug_c_c), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12) 
//

module \ClockDividerP(factor=12)  (bclk, debug_c_c, GND_net) /* synthesis syn_module_defined=1 */ ;
    output bclk;
    input debug_c_c;
    input GND_net;
    
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n50, n40, n54, n48, n36, n7260, n24571;
    wire [31:0]n102;
    
    wire n24570, n24569, n24568, n24567, n24566, n24565, n24564, 
        n24563, n24562, n24561, n24560, n24559, n24558, n24557, 
        n24556, n24184, n24183, n24182, n24181, n24180, n14360, 
        n24179, n24178, n24177, n24176, n24175, n24174, n24173, 
        n24172, n24171, n24170, n24169, n55, n56, n4, n52, n44, 
        n35, n46, n32;
    
    LUT4 i25_4_lut (.A(count[25]), .B(n50), .C(n40), .D(count[9]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(count[7]), .B(count[19]), .C(count[11]), .D(count[21]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[8]), .B(count[29]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i21_4_lut (.A(count[2]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i11_2_lut (.A(count[10]), .B(count[17]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i11_2_lut.init = 16'heeee;
    FD1S3AX clk_o_14 (.D(n7260), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D count_2173_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24571), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_33.INIT1 = 16'h0000;
    defparam count_2173_add_4_33.INJECT1_0 = "NO";
    defparam count_2173_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24570), .COUT(n24571), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2173_add_4_31.INJECT1_0 = "NO";
    defparam count_2173_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24569), .COUT(n24570), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2173_add_4_29.INJECT1_0 = "NO";
    defparam count_2173_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24568), .COUT(n24569), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2173_add_4_27.INJECT1_0 = "NO";
    defparam count_2173_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24567), .COUT(n24568), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2173_add_4_25.INJECT1_0 = "NO";
    defparam count_2173_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24566), .COUT(n24567), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2173_add_4_23.INJECT1_0 = "NO";
    defparam count_2173_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24565), .COUT(n24566), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2173_add_4_21.INJECT1_0 = "NO";
    defparam count_2173_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24564), .COUT(n24565), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2173_add_4_19.INJECT1_0 = "NO";
    defparam count_2173_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24563), .COUT(n24564), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2173_add_4_17.INJECT1_0 = "NO";
    defparam count_2173_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24562), .COUT(n24563), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2173_add_4_15.INJECT1_0 = "NO";
    defparam count_2173_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24561), .COUT(n24562), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2173_add_4_13.INJECT1_0 = "NO";
    defparam count_2173_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24560), .COUT(n24561), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2173_add_4_11.INJECT1_0 = "NO";
    defparam count_2173_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24559), .COUT(n24560), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2173_add_4_9.INJECT1_0 = "NO";
    defparam count_2173_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24558), .COUT(n24559), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2173_add_4_7.INJECT1_0 = "NO";
    defparam count_2173_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24557), .COUT(n24558), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2173_add_4_5.INJECT1_0 = "NO";
    defparam count_2173_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24556), .COUT(n24557), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2173_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2173_add_4_3.INJECT1_0 = "NO";
    defparam count_2173_add_4_3.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24184), .S0(n7260));
    defparam sub_1732_add_2_cout.INIT0 = 16'h0000;
    defparam sub_1732_add_2_cout.INIT1 = 16'h0000;
    defparam sub_1732_add_2_cout.INJECT1_0 = "NO";
    defparam sub_1732_add_2_cout.INJECT1_1 = "NO";
    CCU2D count_2173_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24556), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173_add_4_1.INIT0 = 16'hF000;
    defparam count_2173_add_4_1.INIT1 = 16'h0555;
    defparam count_2173_add_4_1.INJECT1_0 = "NO";
    defparam count_2173_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24183), .COUT(n24184));
    defparam sub_1732_add_2_32.INIT0 = 16'h5555;
    defparam sub_1732_add_2_32.INIT1 = 16'h5555;
    defparam sub_1732_add_2_32.INJECT1_0 = "NO";
    defparam sub_1732_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24182), .COUT(n24183));
    defparam sub_1732_add_2_30.INIT0 = 16'h5555;
    defparam sub_1732_add_2_30.INIT1 = 16'h5555;
    defparam sub_1732_add_2_30.INJECT1_0 = "NO";
    defparam sub_1732_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24181), .COUT(n24182));
    defparam sub_1732_add_2_28.INIT0 = 16'h5555;
    defparam sub_1732_add_2_28.INIT1 = 16'h5555;
    defparam sub_1732_add_2_28.INJECT1_0 = "NO";
    defparam sub_1732_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24180), .COUT(n24181));
    defparam sub_1732_add_2_26.INIT0 = 16'h5555;
    defparam sub_1732_add_2_26.INIT1 = 16'h5555;
    defparam sub_1732_add_2_26.INJECT1_0 = "NO";
    defparam sub_1732_add_2_26.INJECT1_1 = "NO";
    FD1S3IX count_2173__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i1.GSR = "ENABLED";
    CCU2D sub_1732_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24179), .COUT(n24180));
    defparam sub_1732_add_2_24.INIT0 = 16'h5555;
    defparam sub_1732_add_2_24.INIT1 = 16'h5555;
    defparam sub_1732_add_2_24.INJECT1_0 = "NO";
    defparam sub_1732_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24178), .COUT(n24179));
    defparam sub_1732_add_2_22.INIT0 = 16'h5555;
    defparam sub_1732_add_2_22.INIT1 = 16'h5555;
    defparam sub_1732_add_2_22.INJECT1_0 = "NO";
    defparam sub_1732_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24177), .COUT(n24178));
    defparam sub_1732_add_2_20.INIT0 = 16'h5555;
    defparam sub_1732_add_2_20.INIT1 = 16'h5555;
    defparam sub_1732_add_2_20.INJECT1_0 = "NO";
    defparam sub_1732_add_2_20.INJECT1_1 = "NO";
    FD1S3IX count_2173__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i2.GSR = "ENABLED";
    FD1S3IX count_2173__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i3.GSR = "ENABLED";
    FD1S3IX count_2173__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i4.GSR = "ENABLED";
    FD1S3IX count_2173__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i5.GSR = "ENABLED";
    FD1S3IX count_2173__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i6.GSR = "ENABLED";
    FD1S3IX count_2173__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i7.GSR = "ENABLED";
    FD1S3IX count_2173__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i8.GSR = "ENABLED";
    FD1S3IX count_2173__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i9.GSR = "ENABLED";
    FD1S3IX count_2173__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i10.GSR = "ENABLED";
    FD1S3IX count_2173__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i11.GSR = "ENABLED";
    FD1S3IX count_2173__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i12.GSR = "ENABLED";
    FD1S3IX count_2173__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i13.GSR = "ENABLED";
    FD1S3IX count_2173__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i14.GSR = "ENABLED";
    FD1S3IX count_2173__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i15.GSR = "ENABLED";
    FD1S3IX count_2173__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i16.GSR = "ENABLED";
    FD1S3IX count_2173__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i17.GSR = "ENABLED";
    FD1S3IX count_2173__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i18.GSR = "ENABLED";
    FD1S3IX count_2173__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i19.GSR = "ENABLED";
    FD1S3IX count_2173__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i20.GSR = "ENABLED";
    FD1S3IX count_2173__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i21.GSR = "ENABLED";
    FD1S3IX count_2173__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i22.GSR = "ENABLED";
    FD1S3IX count_2173__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i23.GSR = "ENABLED";
    FD1S3IX count_2173__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i24.GSR = "ENABLED";
    FD1S3IX count_2173__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i25.GSR = "ENABLED";
    FD1S3IX count_2173__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i26.GSR = "ENABLED";
    FD1S3IX count_2173__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i27.GSR = "ENABLED";
    FD1S3IX count_2173__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i28.GSR = "ENABLED";
    FD1S3IX count_2173__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i29.GSR = "ENABLED";
    FD1S3IX count_2173__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i30.GSR = "ENABLED";
    FD1S3IX count_2173__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i31.GSR = "ENABLED";
    CCU2D sub_1732_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24176), .COUT(n24177));
    defparam sub_1732_add_2_18.INIT0 = 16'h5555;
    defparam sub_1732_add_2_18.INIT1 = 16'h5555;
    defparam sub_1732_add_2_18.INJECT1_0 = "NO";
    defparam sub_1732_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24175), .COUT(n24176));
    defparam sub_1732_add_2_16.INIT0 = 16'h5555;
    defparam sub_1732_add_2_16.INIT1 = 16'h5555;
    defparam sub_1732_add_2_16.INJECT1_0 = "NO";
    defparam sub_1732_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24174), .COUT(n24175));
    defparam sub_1732_add_2_14.INIT0 = 16'h5555;
    defparam sub_1732_add_2_14.INIT1 = 16'h5555;
    defparam sub_1732_add_2_14.INJECT1_0 = "NO";
    defparam sub_1732_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24173), .COUT(n24174));
    defparam sub_1732_add_2_12.INIT0 = 16'h5555;
    defparam sub_1732_add_2_12.INIT1 = 16'h5555;
    defparam sub_1732_add_2_12.INJECT1_0 = "NO";
    defparam sub_1732_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24172), .COUT(n24173));
    defparam sub_1732_add_2_10.INIT0 = 16'h5555;
    defparam sub_1732_add_2_10.INIT1 = 16'h5555;
    defparam sub_1732_add_2_10.INJECT1_0 = "NO";
    defparam sub_1732_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24171), .COUT(n24172));
    defparam sub_1732_add_2_8.INIT0 = 16'h5555;
    defparam sub_1732_add_2_8.INIT1 = 16'h5555;
    defparam sub_1732_add_2_8.INJECT1_0 = "NO";
    defparam sub_1732_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24170), .COUT(n24171));
    defparam sub_1732_add_2_6.INIT0 = 16'h5555;
    defparam sub_1732_add_2_6.INIT1 = 16'h5555;
    defparam sub_1732_add_2_6.INJECT1_0 = "NO";
    defparam sub_1732_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24169), .COUT(n24170));
    defparam sub_1732_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_1732_add_2_4.INIT1 = 16'h5555;
    defparam sub_1732_add_2_4.INJECT1_0 = "NO";
    defparam sub_1732_add_2_4.INJECT1_1 = "NO";
    FD1S3IX count_2173__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n14360), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2173__i0.GSR = "ENABLED";
    CCU2D sub_1732_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24169));
    defparam sub_1732_add_2_2.INIT0 = 16'h0000;
    defparam sub_1732_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_1732_add_2_2.INJECT1_0 = "NO";
    defparam sub_1732_add_2_2.INJECT1_1 = "NO";
    LUT4 i21306_4_lut (.A(n55), .B(count[1]), .C(n56), .D(n4), .Z(n14360)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i21306_4_lut.init = 16'h0400;
    LUT4 i26_4_lut (.A(count[14]), .B(n52), .C(n44), .D(count[6]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i27_4_lut (.A(n35), .B(n54), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(count[3]), .B(count[0]), .Z(n4)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i23_4_lut (.A(count[24]), .B(n46), .C(n32), .D(count[16]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i15_3_lut (.A(count[15]), .B(count[31]), .C(count[5]), .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i17_4_lut (.A(count[26]), .B(count[12]), .C(count[28]), .D(count[18]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[13]), .B(count[22]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(count[20]), .B(count[4]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i6_2_lut.init = 16'heeee;
    
endmodule
//
// Verilog Description of module \UARTReceiver(baud_div=12) 
//

module \UARTReceiver(baud_div=12)  (debug_c_7, n1315, n1316, n10741, 
            n9388_c, debug_c_c, n28981, rx_data, n28952, n30646, 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    output debug_c_7;
    input n1315;
    input n1316;
    output n10741;
    input n9388_c;
    input debug_c_c;
    input n28981;
    output [7:0]rx_data;
    input n28952;
    input n30646;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n25707, n13501;
    wire [5:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    
    wire n13502, n32, bclk, n27992;
    wire [7:0]rdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(22[12:17])
    
    wire n27993, n54;
    wire [7:0]n78;
    
    wire n11674, n13, n7926, n29045, n29050, n28988;
    wire [5:0]n23;
    
    wire n29, n29030, n29001, n28547, n28546, n28887, n7928, n25915, 
        baud_reset, n86_adj_268, n18, n20, n13881, n25847, n27981, 
        n7968, n7966, n7964, n7962, n7960, n7958, n7956, n7954, 
        n7952, n7950, n7948, n7946, n7944, n7942, n29044, n27307, 
        n27085, n27979, n27980, n11683, n19, n88, n28980, n55, 
        n24725, n56, n2683;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n52, n44, n35, n54_adj_269, n48, n36, n46, n32_adj_270, 
        n50, n40, n26345, n13880;
    
    PFUMX i7736 (.BLUT(n25707), .ALUT(n13501), .C0(state[0]), .Z(n13502));
    LUT4 i1_4_lut (.A(state[4]), .B(state[3]), .C(state[2]), .D(state[1]), 
         .Z(n32)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut.init = 16'heaaa;
    LUT4 rdata_1__bdd_3_lut_4_lut (.A(state[1]), .B(bclk), .C(n27992), 
         .D(rdata[1]), .Z(n27993)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam rdata_1__bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut (.A(state[1]), .B(bclk), .C(state[2]), .Z(n54)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_3_lut (.A(debug_c_7), .B(n1315), .C(n1316), .Z(n10741)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_3_lut.init = 16'h5454;
    LUT4 i1_4_lut_adj_263 (.A(n78[0]), .B(rdata[0]), .C(n11674), .D(n13), 
         .Z(n7926)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_263.init = 16'heca0;
    LUT4 i3818_4_lut (.A(n9388_c), .B(rdata[0]), .C(n29045), .D(n29050), 
         .Z(n78[0])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3818_4_lut.init = 16'hccca;
    LUT4 i2_3_lut (.A(state[5]), .B(state[4]), .C(state[0]), .Z(n11674)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i2_3_lut.init = 16'h0404;
    LUT4 i2_3_lut_adj_264 (.A(state[0]), .B(state[5]), .C(state[4]), .Z(n13)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_3_lut_adj_264.init = 16'hefef;
    LUT4 i18248_4_lut (.A(n28988), .B(state[5]), .C(n23[3]), .D(n32), 
         .Z(n29)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i18248_4_lut.init = 16'h3111;
    LUT4 i2919_3_lut_rep_372 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n29030)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2919_3_lut_rep_372.init = 16'h8080;
    LUT4 i2926_2_lut_rep_343_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(state[3]), .Z(n29001)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2926_2_lut_rep_343_4_lut.init = 16'h8000;
    FD1P3AX rdata_i0_i0 (.D(n7926), .SP(n28981), .CK(debug_c_c), .Q(rdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i0.GSR = "ENABLED";
    LUT4 n28547_bdd_4_lut (.A(n28547), .B(n32), .C(n28546), .D(state[0]), 
         .Z(n28887)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;
    defparam n28547_bdd_4_lut.init = 16'hf088;
    FD1P3AX data_i0_i0 (.D(n7928), .SP(n28981), .CK(debug_c_c), .Q(rx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i0.GSR = "ENABLED";
    FD1S3IX state__i0 (.D(n25915), .CK(debug_c_c), .CD(n28952), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i0.GSR = "ENABLED";
    FD1S3JX baud_reset_52 (.D(n86_adj_268), .CK(debug_c_c), .PD(n28952), 
            .Q(baud_reset)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam baud_reset_52.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_265 (.A(state[5]), .B(state[2]), .C(n28988), .D(n32), 
         .Z(n18)) /* synthesis lut_function=(!(A+!(B ((D)+!C)+!B !(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_265.init = 16'h4505;
    LUT4 i33_3_lut (.A(state[1]), .B(state[2]), .C(bclk), .Z(n20)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i33_3_lut.init = 16'hc6c6;
    FD1S3IX state__i5 (.D(n13502), .CK(debug_c_c), .CD(n28952), .Q(state[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i5.GSR = "ENABLED";
    FD1S3IX state__i4 (.D(n28887), .CK(debug_c_c), .CD(n28952), .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i4.GSR = "ENABLED";
    FD1S3IX state__i3 (.D(n13881), .CK(debug_c_c), .CD(n28952), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i3.GSR = "ENABLED";
    FD1S3IX state__i2 (.D(n25847), .CK(debug_c_c), .CD(n30646), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i2.GSR = "ENABLED";
    FD1S3IX state__i1 (.D(n27981), .CK(debug_c_c), .CD(n30646), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i1.GSR = "ENABLED";
    FD1P3AX data_i0_i7 (.D(n7968), .SP(n28981), .CK(debug_c_c), .Q(rx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i7.GSR = "ENABLED";
    FD1P3AX data_i0_i6 (.D(n7966), .SP(n28981), .CK(debug_c_c), .Q(rx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i6.GSR = "ENABLED";
    FD1P3AX data_i0_i5 (.D(n7964), .SP(n28981), .CK(debug_c_c), .Q(rx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i5.GSR = "ENABLED";
    FD1P3AX data_i0_i4 (.D(n7962), .SP(n28981), .CK(debug_c_c), .Q(rx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i4.GSR = "ENABLED";
    FD1P3AX data_i0_i3 (.D(n7960), .SP(n28981), .CK(debug_c_c), .Q(rx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i3.GSR = "ENABLED";
    FD1P3AX data_i0_i2 (.D(n7958), .SP(n28981), .CK(debug_c_c), .Q(rx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i2.GSR = "ENABLED";
    FD1P3AX data_i0_i1 (.D(n7956), .SP(n28981), .CK(debug_c_c), .Q(rx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i1.GSR = "ENABLED";
    FD1P3AX rdata_i0_i7 (.D(n7954), .SP(n28981), .CK(debug_c_c), .Q(rdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i7.GSR = "ENABLED";
    FD1P3AX rdata_i0_i6 (.D(n7952), .SP(n28981), .CK(debug_c_c), .Q(rdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i6.GSR = "ENABLED";
    FD1P3AX rdata_i0_i5 (.D(n7950), .SP(n28981), .CK(debug_c_c), .Q(rdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i5.GSR = "ENABLED";
    FD1P3AX rdata_i0_i4 (.D(n7948), .SP(n28981), .CK(debug_c_c), .Q(rdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i4.GSR = "ENABLED";
    FD1P3AX rdata_i0_i3 (.D(n7946), .SP(n28981), .CK(debug_c_c), .Q(rdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i3.GSR = "ENABLED";
    FD1P3AX rdata_i0_i2 (.D(n7944), .SP(n28981), .CK(debug_c_c), .Q(rdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i2.GSR = "ENABLED";
    FD1P3AX rdata_i0_i1 (.D(n7942), .SP(n28981), .CK(debug_c_c), .Q(rdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_386 (.A(state[1]), .B(state[4]), .Z(n29044)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_rep_386.init = 16'heeee;
    LUT4 i1_2_lut_rep_330_3_lut_4_lut (.A(state[1]), .B(state[4]), .C(n9388_c), 
         .D(n29045), .Z(n28988)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_rep_330_3_lut_4_lut.init = 16'hfffe;
    LUT4 i20937_3_lut_4_lut (.A(state[1]), .B(state[4]), .C(n29045), .D(n9388_c), 
         .Z(n27307)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i20937_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_387 (.A(state[2]), .B(state[3]), .Z(n29045)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_rep_387.init = 16'heeee;
    LUT4 i1_2_lut_rep_392 (.A(state[1]), .B(bclk), .Z(n29050)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i1_2_lut_rep_392.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_adj_266 (.A(state[1]), .B(bclk), .C(state[2]), 
         .Z(n27085)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i1_2_lut_3_lut_adj_266.init = 16'hbfbf;
    LUT4 n116_bdd_2_lut (.A(state[1]), .B(bclk), .Z(n27979)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam n116_bdd_2_lut.init = 16'h9999;
    LUT4 n116_bdd_4_lut_21682 (.A(n28988), .B(state[1]), .C(n32), .D(state[5]), 
         .Z(n27980)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (D))) */ ;
    defparam n116_bdd_4_lut_21682.init = 16'h00d5;
    LUT4 i1_4_lut_adj_267 (.A(rdata[0]), .B(rx_data[0]), .C(n11683), .D(n19), 
         .Z(n7928)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_267.init = 16'heca0;
    LUT4 i4_4_lut (.A(n29045), .B(n29044), .C(state[5]), .D(state[0]), 
         .Z(n19)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i4_4_lut.init = 16'hffef;
    LUT4 i1_4_lut_adj_268 (.A(bclk), .B(state[0]), .C(state[5]), .D(n32), 
         .Z(n25915)) /* synthesis lut_function=(A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_268.init = 16'h8a88;
    LUT4 i1_4_lut_adj_269 (.A(rdata[7]), .B(rx_data[7]), .C(n11683), .D(n19), 
         .Z(n7968)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_269.init = 16'heca0;
    LUT4 i1_4_lut_adj_270 (.A(rdata[6]), .B(rx_data[6]), .C(n11683), .D(n19), 
         .Z(n7966)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_270.init = 16'heca0;
    LUT4 i1_4_lut_adj_271 (.A(rdata[5]), .B(rx_data[5]), .C(n11683), .D(n19), 
         .Z(n7964)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_271.init = 16'heca0;
    LUT4 i1_4_lut_adj_272 (.A(rdata[4]), .B(rx_data[4]), .C(n11683), .D(n19), 
         .Z(n7962)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_272.init = 16'heca0;
    LUT4 i1_4_lut_adj_273 (.A(rdata[3]), .B(rx_data[3]), .C(n11683), .D(n19), 
         .Z(n7960)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_273.init = 16'heca0;
    LUT4 i1_4_lut_adj_274 (.A(rdata[2]), .B(rx_data[2]), .C(n11683), .D(n19), 
         .Z(n7958)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_274.init = 16'heca0;
    LUT4 i1_4_lut_adj_275 (.A(rdata[1]), .B(rx_data[1]), .C(n11683), .D(n19), 
         .Z(n7956)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_275.init = 16'heca0;
    FD1S3IX drdy_51 (.D(n88), .CK(debug_c_c), .CD(n30646), .Q(debug_c_7));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam drdy_51.GSR = "ENABLED";
    LUT4 n113_bdd_4_lut (.A(n9388_c), .B(state[2]), .C(rdata[1]), .D(state[3]), 
         .Z(n27992)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)))) */ ;
    defparam n113_bdd_4_lut.init = 16'hf0e2;
    LUT4 i7735_3_lut_4_lut (.A(state[4]), .B(n29001), .C(bclk), .D(state[5]), 
         .Z(n13501)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;
    defparam i7735_3_lut_4_lut.init = 16'hf708;
    LUT4 i21183_4_lut (.A(bclk), .B(n27307), .C(state[5]), .D(n28980), 
         .Z(n25707)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i21183_4_lut.init = 16'h3a30;
    LUT4 i1_4_lut_adj_276 (.A(baud_reset), .B(n55), .C(n24725), .D(n56), 
         .Z(n2683)) /* synthesis lut_function=(A+!(B+((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_276.init = 16'haaba;
    LUT4 i1_4_lut_adj_277 (.A(n78[7]), .B(rdata[7]), .C(n11674), .D(n13), 
         .Z(n7954)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_277.init = 16'heca0;
    LUT4 i26_4_lut (.A(count[2]), .B(n52), .C(n44), .D(count[15]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i3679_4_lut (.A(rdata[7]), .B(n9388_c), .C(state[3]), .D(n54), 
         .Z(n78[7])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3679_4_lut.init = 16'hcaaa;
    LUT4 i27_4_lut (.A(n35), .B(n54_adj_269), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i23_4_lut (.A(count[13]), .B(n46), .C(n32_adj_270), .D(count[22]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i15_3_lut (.A(count[6]), .B(count[5]), .C(count[31]), .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i17_4_lut (.A(count[24]), .B(count[29]), .C(count[16]), .D(count[7]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[26]), .B(count[28]), .Z(n32_adj_270)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_278 (.A(n78[6]), .B(rdata[6]), .C(n11674), .D(n13), 
         .Z(n7952)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_278.init = 16'heca0;
    LUT4 i6_2_lut (.A(count[11]), .B(count[19]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i25_4_lut (.A(count[8]), .B(n50), .C(n40), .D(count[23]), .Z(n54_adj_269)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(count[12]), .B(count[20]), .C(count[18]), .D(count[4]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[21]), .B(count[25]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i21_4_lut (.A(count[14]), .B(count[10]), .C(count[9]), .D(count[17]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i3681_4_lut (.A(n9388_c), .B(rdata[6]), .C(state[3]), .D(n27085), 
         .Z(n78[6])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3681_4_lut.init = 16'hccac;
    LUT4 i11_2_lut (.A(count[27]), .B(count[30]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i11_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_279 (.A(n78[5]), .B(rdata[5]), .C(n11674), .D(n13), 
         .Z(n7950)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_279.init = 16'heca0;
    LUT4 i3683_4_lut (.A(n9388_c), .B(rdata[5]), .C(state[1]), .D(n26345), 
         .Z(n78[5])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3683_4_lut.init = 16'hccac;
    LUT4 i2_3_lut_adj_280 (.A(bclk), .B(state[3]), .C(state[2]), .Z(n26345)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i2_3_lut_adj_280.init = 16'hf7f7;
    LUT4 i1_4_lut_adj_281 (.A(n78[4]), .B(rdata[4]), .C(n11674), .D(n13), 
         .Z(n7948)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_281.init = 16'heca0;
    LUT4 i3685_4_lut (.A(n9388_c), .B(rdata[4]), .C(state[1]), .D(n26345), 
         .Z(n78[4])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3685_4_lut.init = 16'hccca;
    LUT4 i1_4_lut_adj_282 (.A(n78[3]), .B(rdata[3]), .C(n11674), .D(n13), 
         .Z(n7946)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_282.init = 16'heca0;
    LUT4 i3687_4_lut (.A(n9388_c), .B(rdata[3]), .C(state[3]), .D(n54), 
         .Z(n78[3])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3687_4_lut.init = 16'hcacc;
    LUT4 i1_4_lut_adj_283 (.A(n78[2]), .B(rdata[2]), .C(n11674), .D(n13), 
         .Z(n7944)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_283.init = 16'heca0;
    LUT4 i3689_4_lut (.A(n9388_c), .B(rdata[2]), .C(state[3]), .D(n27085), 
         .Z(n78[2])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3689_4_lut.init = 16'hccca;
    LUT4 i1_4_lut_adj_284 (.A(n27993), .B(rdata[1]), .C(n11674), .D(n13), 
         .Z(n7942)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_284.init = 16'heca0;
    LUT4 n32_bdd_3_lut_21717_4_lut (.A(state[3]), .B(n29030), .C(bclk), 
         .D(state[4]), .Z(n28546)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;
    defparam n32_bdd_3_lut_21717_4_lut.init = 16'hf708;
    LUT4 i2933_2_lut_rep_322_3_lut (.A(state[3]), .B(n29030), .C(state[4]), 
         .Z(n28980)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2933_2_lut_rep_322_3_lut.init = 16'h8080;
    LUT4 i2_3_lut_4_lut (.A(n29045), .B(n29044), .C(state[0]), .D(state[5]), 
         .Z(n11683)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i2_3_lut_4_lut.init = 16'h0100;
    LUT4 mux_8_i4_3_lut_3_lut (.A(state[3]), .B(n29030), .C(bclk), .Z(n23[3])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;
    defparam mux_8_i4_3_lut_3_lut.init = 16'h6a6a;
    LUT4 i8114_3_lut_3_lut (.A(state[3]), .B(n29030), .C(bclk), .Z(n13880)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;
    defparam i8114_3_lut_3_lut.init = 16'ha6a6;
    PFUMX i8115 (.BLUT(n29), .ALUT(n13880), .C0(state[0]), .Z(n13881));
    PFUMX i32 (.BLUT(n18), .ALUT(n20), .C0(state[0]), .Z(n25847));
    LUT4 n32_bdd_4_lut_21718 (.A(state[4]), .B(state[5]), .C(bclk), .D(n29001), 
         .Z(n28547)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+!(C (D))))) */ ;
    defparam n32_bdd_4_lut_21718.init = 16'h1222;
    LUT4 i1_3_lut_4_lut (.A(state[0]), .B(n28988), .C(baud_reset), .D(n11683), 
         .Z(n86_adj_268)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[13:20])
    defparam i1_3_lut_4_lut.init = 16'hffe0;
    LUT4 i1_3_lut_4_lut_adj_285 (.A(state[0]), .B(n28988), .C(debug_c_7), 
         .D(n11683), .Z(n88)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[13:20])
    defparam i1_3_lut_4_lut_adj_285.init = 16'hffe0;
    PFUMX i21468 (.BLUT(n27980), .ALUT(n27979), .C0(state[0]), .Z(n27981));
    \ClockDividerP(factor=12)_U0  baud_gen (.count({count[31:5], Open_59, 
            Open_60, Open_61, Open_62, Open_63}), .GND_net(GND_net), 
            .\count[4] (count[4]), .\count[2] (count[2]), .bclk(bclk), 
            .debug_c_c(debug_c_c), .baud_reset(baud_reset), .n24725(n24725), 
            .n2683(n2683)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(25[28] 27[56])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12)_U0 
//

module \ClockDividerP(factor=12)_U0  (count, GND_net, \count[4] , \count[2] , 
            bclk, debug_c_c, baud_reset, n24725, n2683) /* synthesis syn_module_defined=1 */ ;
    output [31:0]count;
    input GND_net;
    output \count[4] ;
    output \count[2] ;
    output bclk;
    input debug_c_c;
    input baud_reset;
    output n24725;
    input n2683;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n24523;
    wire [31:0]n134;
    
    wire n24522, n24521, n24520, n24519, n24518, n24517, n24516, 
        n24515, n24514, n24513, n24512, n24511, n24510, n24509;
    wire [31:0]count_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n24508, n7225, n24200, n24199, n24198, n24197, n24196, 
        n24195, n24194, n24193, n24192, n24191, n24190, n24189, 
        n24188, n24187, n24186, n24185;
    
    CCU2D count_2172_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24523), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_33.INIT1 = 16'h0000;
    defparam count_2172_add_4_33.INJECT1_0 = "NO";
    defparam count_2172_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24522), .COUT(n24523), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2172_add_4_31.INJECT1_0 = "NO";
    defparam count_2172_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24521), .COUT(n24522), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2172_add_4_29.INJECT1_0 = "NO";
    defparam count_2172_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24520), .COUT(n24521), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2172_add_4_27.INJECT1_0 = "NO";
    defparam count_2172_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24519), .COUT(n24520), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2172_add_4_25.INJECT1_0 = "NO";
    defparam count_2172_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24518), .COUT(n24519), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2172_add_4_23.INJECT1_0 = "NO";
    defparam count_2172_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24517), .COUT(n24518), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2172_add_4_21.INJECT1_0 = "NO";
    defparam count_2172_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24516), .COUT(n24517), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2172_add_4_19.INJECT1_0 = "NO";
    defparam count_2172_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24515), .COUT(n24516), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2172_add_4_17.INJECT1_0 = "NO";
    defparam count_2172_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24514), .COUT(n24515), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2172_add_4_15.INJECT1_0 = "NO";
    defparam count_2172_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24513), .COUT(n24514), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2172_add_4_13.INJECT1_0 = "NO";
    defparam count_2172_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24512), .COUT(n24513), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2172_add_4_11.INJECT1_0 = "NO";
    defparam count_2172_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24511), .COUT(n24512), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2172_add_4_9.INJECT1_0 = "NO";
    defparam count_2172_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24510), .COUT(n24511), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2172_add_4_7.INJECT1_0 = "NO";
    defparam count_2172_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_5 (.A0(count_c[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count[4] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24509), .COUT(n24510), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2172_add_4_5.INJECT1_0 = "NO";
    defparam count_2172_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_3 (.A0(count_c[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count[2] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24508), .COUT(n24509), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2172_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2172_add_4_3.INJECT1_0 = "NO";
    defparam count_2172_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2172_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n24508), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172_add_4_1.INIT0 = 16'hF000;
    defparam count_2172_add_4_1.INIT1 = 16'h0555;
    defparam count_2172_add_4_1.INJECT1_0 = "NO";
    defparam count_2172_add_4_1.INJECT1_1 = "NO";
    FD1S3IX clk_o_14 (.D(n7225), .CK(debug_c_c), .CD(baud_reset), .Q(bclk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    LUT4 i2_3_lut (.A(count_c[1]), .B(count_c[3]), .C(count_c[0]), .Z(n24725)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    FD1S3IX count_2172__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2683), .Q(count_c[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i0.GSR = "ENABLED";
    CCU2D sub_1730_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24200), .S0(n7225));
    defparam sub_1730_add_2_cout.INIT0 = 16'h0000;
    defparam sub_1730_add_2_cout.INIT1 = 16'h0000;
    defparam sub_1730_add_2_cout.INJECT1_0 = "NO";
    defparam sub_1730_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_1730_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24199), .COUT(n24200));
    defparam sub_1730_add_2_32.INIT0 = 16'h5555;
    defparam sub_1730_add_2_32.INIT1 = 16'h5555;
    defparam sub_1730_add_2_32.INJECT1_0 = "NO";
    defparam sub_1730_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_1730_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24198), .COUT(n24199));
    defparam sub_1730_add_2_30.INIT0 = 16'h5555;
    defparam sub_1730_add_2_30.INIT1 = 16'h5555;
    defparam sub_1730_add_2_30.INJECT1_0 = "NO";
    defparam sub_1730_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_1730_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24197), .COUT(n24198));
    defparam sub_1730_add_2_28.INIT0 = 16'h5555;
    defparam sub_1730_add_2_28.INIT1 = 16'h5555;
    defparam sub_1730_add_2_28.INJECT1_0 = "NO";
    defparam sub_1730_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_1730_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24196), .COUT(n24197));
    defparam sub_1730_add_2_26.INIT0 = 16'h5555;
    defparam sub_1730_add_2_26.INIT1 = 16'h5555;
    defparam sub_1730_add_2_26.INJECT1_0 = "NO";
    defparam sub_1730_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_1730_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24195), .COUT(n24196));
    defparam sub_1730_add_2_24.INIT0 = 16'h5555;
    defparam sub_1730_add_2_24.INIT1 = 16'h5555;
    defparam sub_1730_add_2_24.INJECT1_0 = "NO";
    defparam sub_1730_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_1730_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24194), .COUT(n24195));
    defparam sub_1730_add_2_22.INIT0 = 16'h5555;
    defparam sub_1730_add_2_22.INIT1 = 16'h5555;
    defparam sub_1730_add_2_22.INJECT1_0 = "NO";
    defparam sub_1730_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_1730_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24193), .COUT(n24194));
    defparam sub_1730_add_2_20.INIT0 = 16'h5555;
    defparam sub_1730_add_2_20.INIT1 = 16'h5555;
    defparam sub_1730_add_2_20.INJECT1_0 = "NO";
    defparam sub_1730_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_1730_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24192), .COUT(n24193));
    defparam sub_1730_add_2_18.INIT0 = 16'h5555;
    defparam sub_1730_add_2_18.INIT1 = 16'h5555;
    defparam sub_1730_add_2_18.INJECT1_0 = "NO";
    defparam sub_1730_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_1730_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24191), .COUT(n24192));
    defparam sub_1730_add_2_16.INIT0 = 16'h5555;
    defparam sub_1730_add_2_16.INIT1 = 16'h5555;
    defparam sub_1730_add_2_16.INJECT1_0 = "NO";
    defparam sub_1730_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_1730_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24190), .COUT(n24191));
    defparam sub_1730_add_2_14.INIT0 = 16'h5555;
    defparam sub_1730_add_2_14.INIT1 = 16'h5555;
    defparam sub_1730_add_2_14.INJECT1_0 = "NO";
    defparam sub_1730_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_1730_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24189), .COUT(n24190));
    defparam sub_1730_add_2_12.INIT0 = 16'h5555;
    defparam sub_1730_add_2_12.INIT1 = 16'h5555;
    defparam sub_1730_add_2_12.INJECT1_0 = "NO";
    defparam sub_1730_add_2_12.INJECT1_1 = "NO";
    FD1S3IX count_2172__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2683), .Q(count_c[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i1.GSR = "ENABLED";
    CCU2D sub_1730_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24188), .COUT(n24189));
    defparam sub_1730_add_2_10.INIT0 = 16'h5555;
    defparam sub_1730_add_2_10.INIT1 = 16'h5555;
    defparam sub_1730_add_2_10.INJECT1_0 = "NO";
    defparam sub_1730_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_1730_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24187), .COUT(n24188));
    defparam sub_1730_add_2_8.INIT0 = 16'h5555;
    defparam sub_1730_add_2_8.INIT1 = 16'h5555;
    defparam sub_1730_add_2_8.INJECT1_0 = "NO";
    defparam sub_1730_add_2_8.INJECT1_1 = "NO";
    FD1S3IX count_2172__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2683), .Q(\count[2] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i2.GSR = "ENABLED";
    FD1S3IX count_2172__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2683), .Q(count_c[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i3.GSR = "ENABLED";
    FD1S3IX count_2172__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2683), .Q(\count[4] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i4.GSR = "ENABLED";
    FD1S3IX count_2172__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2683), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i5.GSR = "ENABLED";
    FD1S3IX count_2172__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2683), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i6.GSR = "ENABLED";
    FD1S3IX count_2172__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2683), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i7.GSR = "ENABLED";
    FD1S3IX count_2172__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2683), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i8.GSR = "ENABLED";
    FD1S3IX count_2172__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2683), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i9.GSR = "ENABLED";
    FD1S3IX count_2172__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i10.GSR = "ENABLED";
    FD1S3IX count_2172__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i11.GSR = "ENABLED";
    FD1S3IX count_2172__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i12.GSR = "ENABLED";
    FD1S3IX count_2172__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i13.GSR = "ENABLED";
    FD1S3IX count_2172__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i14.GSR = "ENABLED";
    FD1S3IX count_2172__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i15.GSR = "ENABLED";
    FD1S3IX count_2172__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i16.GSR = "ENABLED";
    FD1S3IX count_2172__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i17.GSR = "ENABLED";
    FD1S3IX count_2172__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i18.GSR = "ENABLED";
    FD1S3IX count_2172__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i19.GSR = "ENABLED";
    FD1S3IX count_2172__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i20.GSR = "ENABLED";
    FD1S3IX count_2172__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i21.GSR = "ENABLED";
    FD1S3IX count_2172__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i22.GSR = "ENABLED";
    FD1S3IX count_2172__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i23.GSR = "ENABLED";
    FD1S3IX count_2172__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i24.GSR = "ENABLED";
    FD1S3IX count_2172__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i25.GSR = "ENABLED";
    FD1S3IX count_2172__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i26.GSR = "ENABLED";
    FD1S3IX count_2172__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i27.GSR = "ENABLED";
    FD1S3IX count_2172__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i28.GSR = "ENABLED";
    FD1S3IX count_2172__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i29.GSR = "ENABLED";
    FD1S3IX count_2172__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i30.GSR = "ENABLED";
    FD1S3IX count_2172__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2683), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2172__i31.GSR = "ENABLED";
    CCU2D sub_1730_add_2_6 (.A0(\count[4] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24186), .COUT(n24187));
    defparam sub_1730_add_2_6.INIT0 = 16'h5555;
    defparam sub_1730_add_2_6.INIT1 = 16'h5555;
    defparam sub_1730_add_2_6.INJECT1_0 = "NO";
    defparam sub_1730_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_1730_add_2_4 (.A0(\count[2] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24185), .COUT(n24186));
    defparam sub_1730_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_1730_add_2_4.INIT1 = 16'h5555;
    defparam sub_1730_add_2_4.INJECT1_0 = "NO";
    defparam sub_1730_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_1730_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[1]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n24185));
    defparam sub_1730_add_2_2.INIT0 = 16'h0000;
    defparam sub_1730_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_1730_add_2_2.INJECT1_0 = "NO";
    defparam sub_1730_add_2_2.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module GlobalControlPeripheral
//

module GlobalControlPeripheral (\select[1] , n30644, n29028, rw, n6, 
            \read_value[2] , debug_c_c, n12042, n8040, read_size, 
            n88, n30649, signal_light_c, n10501, n14439, \control_reg[7] , 
            n24911, stepping, \control_reg[7]_adj_144 , n24994, n21, 
            \control_reg[7]_adj_145 , n24970, stepping_adj_146, n10489, 
            n14286, \control_reg[7]_adj_147 , n24974, stepping_adj_148, 
            \register[2][31] , n30648, \register[2][30] , \register[2][29] , 
            \register[2][28] , \register[2][27] , \register[2][26] , \register[2][25] , 
            \register[2][24] , \register[2][23] , \register[2][22] , \register[2][21] , 
            \register[2][20] , \register[2][19] , \register[2][18] , \register[2][17] , 
            \register[2][16] , \register[2][15] , \register[2][14] , \register[2][13] , 
            \register[2][12] , \register[2][11] , \register[2][10] , \register[2][9] , 
            \register[2][8] , \register[2][7] , \register[2][6] , \register[2][5] , 
            \register[2][4] , \register_addr[0] , n30647, n28991, xbee_pause_c, 
            \register_addr[5] , n28972, \register_addr[1] , \register_addr[2] , 
            n28920, n22447, GND_net, n28921, n29063, n8044, n29025, 
            n29011, n28901, \read_value[3] , \read_value[4] , n27030, 
            \read_value[5] , n27034, n48, \read_value[6] , n27036, 
            n28990, \read_value[7] , n27028, \read_value[8] , n27046, 
            \read_value[9] , n27042, \read_value[10] , n27045, \read_value[11] , 
            n27026, \read_value[12] , n27025, \read_value[13] , n27027, 
            \read_value[14] , n27029, \read_value[15] , n27038, \read_value[16] , 
            n27031, \read_value[17] , n27033, \read_value[18] , n27023, 
            \read_value[19] , n27041, \read_value[20] , n27047, \read_value[21] , 
            n27048, \read_value[22] , n27040, \read_value[23] , n27039, 
            \read_value[24] , n27035, \read_value[25] , n27050, \read_value[26] , 
            n27024, \read_value[27] , n27049, \read_value[28] , n27044, 
            \read_value[29] , n27032, \read_value[30] , n27037, \read_value[31] , 
            n27043, \read_value[0] , n14380, n27065, n14379, \databus[1] ) /* synthesis syn_module_defined=1 */ ;
    input \select[1] ;
    input n30644;
    output n29028;
    input rw;
    output n6;
    output \read_value[2] ;
    input debug_c_c;
    output n12042;
    input n8040;
    output [2:0]read_size;
    input n88;
    input n30649;
    output signal_light_c;
    input n10501;
    output n14439;
    input \control_reg[7] ;
    input n24911;
    output stepping;
    input \control_reg[7]_adj_144 ;
    input n24994;
    output n21;
    input \control_reg[7]_adj_145 ;
    input n24970;
    output stepping_adj_146;
    input n10489;
    output n14286;
    input \control_reg[7]_adj_147 ;
    input n24974;
    output stepping_adj_148;
    output \register[2][31] ;
    input n30648;
    output \register[2][30] ;
    output \register[2][29] ;
    output \register[2][28] ;
    output \register[2][27] ;
    output \register[2][26] ;
    output \register[2][25] ;
    output \register[2][24] ;
    output \register[2][23] ;
    output \register[2][22] ;
    output \register[2][21] ;
    output \register[2][20] ;
    output \register[2][19] ;
    output \register[2][18] ;
    output \register[2][17] ;
    output \register[2][16] ;
    output \register[2][15] ;
    output \register[2][14] ;
    output \register[2][13] ;
    output \register[2][12] ;
    output \register[2][11] ;
    output \register[2][10] ;
    output \register[2][9] ;
    output \register[2][8] ;
    output \register[2][7] ;
    output \register[2][6] ;
    output \register[2][5] ;
    output \register[2][4] ;
    input \register_addr[0] ;
    input n30647;
    input n28991;
    input xbee_pause_c;
    input \register_addr[5] ;
    input n28972;
    input \register_addr[1] ;
    input \register_addr[2] ;
    output n28920;
    input n22447;
    input GND_net;
    input n28921;
    input n29063;
    output n8044;
    input n29025;
    input n29011;
    output n28901;
    output \read_value[3] ;
    output \read_value[4] ;
    input n27030;
    output \read_value[5] ;
    input n27034;
    input n48;
    output \read_value[6] ;
    input n27036;
    input n28990;
    output \read_value[7] ;
    input n27028;
    output \read_value[8] ;
    input n27046;
    output \read_value[9] ;
    input n27042;
    output \read_value[10] ;
    input n27045;
    output \read_value[11] ;
    input n27026;
    output \read_value[12] ;
    input n27025;
    output \read_value[13] ;
    input n27027;
    output \read_value[14] ;
    input n27029;
    output \read_value[15] ;
    input n27038;
    output \read_value[16] ;
    input n27031;
    output \read_value[17] ;
    input n27033;
    output \read_value[18] ;
    input n27023;
    output \read_value[19] ;
    input n27041;
    output \read_value[20] ;
    input n27047;
    output \read_value[21] ;
    input n27048;
    output \read_value[22] ;
    input n27040;
    output \read_value[23] ;
    input n27039;
    output \read_value[24] ;
    input n27035;
    output \read_value[25] ;
    input n27050;
    output \read_value[26] ;
    input n27024;
    output \read_value[27] ;
    input n27049;
    output \read_value[28] ;
    input n27044;
    output \read_value[29] ;
    input n27032;
    output \read_value[30] ;
    input n27037;
    output \read_value[31] ;
    input n27043;
    output \read_value[0] ;
    input n14380;
    input n27065;
    input n14379;
    input \databus[1] ;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(30[13:23])
    
    wire n28060, n28053;
    wire [31:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    
    wire n7991;
    wire [31:0]n100;
    
    wire prev_clk_1Hz, clk_1Hz;
    wire [31:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    
    wire n178, prev_select, force_pause, n29036, n27213, n25733, 
        n15, n24232, n24231, n24230, n24229, n24228, n24227, n24226, 
        n24225, n24224, n24223, n28058, n28051, n24222, n24221, 
        n24220, n24219, n24218, n24217;
    wire [31:0]n6443;
    
    wire n11839, n25965, n21_adj_267;
    
    LUT4 i14_2_lut_rep_370 (.A(\select[1] ), .B(n30644), .Z(n29028)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(35[19:32])
    defparam i14_2_lut_rep_370.init = 16'h8888;
    LUT4 Select_3616_i6_2_lut_3_lut (.A(\select[1] ), .B(rw), .C(read_value[1]), 
         .Z(n6)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(35[19:32])
    defparam Select_3616_i6_2_lut_3_lut.init = 16'h8080;
    FD1P3AX read_value__i2 (.D(n28060), .SP(n12042), .CK(debug_c_c), .Q(\read_value[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n28053), .SP(n12042), .CD(n8040), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3AX read_size_i0_i0 (.D(n88), .SP(n12042), .CK(debug_c_c), .Q(read_size[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i0.GSR = "ENABLED";
    FD1P3IX uptime_count__i0 (.D(n100[0]), .SP(n7991), .CD(n30649), .CK(debug_c_c), 
            .Q(\register[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i0.GSR = "ENABLED";
    FD1S3AX prev_clk_1Hz_149 (.D(clk_1Hz), .CK(debug_c_c), .Q(prev_clk_1Hz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam prev_clk_1Hz_149.GSR = "ENABLED";
    FD1S3AX xbee_pause_latched_150 (.D(n178), .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam xbee_pause_latched_150.GSR = "ENABLED";
    FD1S3AX prev_select_148 (.D(\select[1] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam prev_select_148.GSR = "ENABLED";
    LUT4 i112_2_lut_rep_378 (.A(\register[0] [2]), .B(force_pause), .Z(n29036)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i112_2_lut_rep_378.init = 16'heeee;
    LUT4 i14026_2_lut_3_lut (.A(\register[0] [2]), .B(force_pause), .C(clk_1Hz), 
         .Z(signal_light_c)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i14026_2_lut_3_lut.init = 16'hfefe;
    LUT4 i8678_2_lut_3_lut (.A(\register[0] [2]), .B(force_pause), .C(n10501), 
         .Z(n14439)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i8678_2_lut_3_lut.init = 16'he0e0;
    LUT4 i2_3_lut_4_lut (.A(\register[0] [2]), .B(force_pause), .C(\control_reg[7] ), 
         .D(n24911), .Z(stepping)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut.init = 16'h1000;
    LUT4 i2_3_lut_4_lut_adj_260 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7]_adj_144 ), .D(n24994), .Z(n21)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_260.init = 16'h1000;
    LUT4 i2_3_lut_4_lut_adj_261 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7]_adj_145 ), .D(n24970), .Z(stepping_adj_146)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_261.init = 16'h1000;
    LUT4 i8646_2_lut_3_lut (.A(\register[0] [2]), .B(force_pause), .C(n10489), 
         .Z(n14286)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i8646_2_lut_3_lut.init = 16'he0e0;
    LUT4 i2_3_lut_4_lut_adj_262 (.A(\register[0] [2]), .B(force_pause), 
         .C(\control_reg[7]_adj_147 ), .D(n24974), .Z(stepping_adj_148)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_262.init = 16'h1000;
    FD1P3IX uptime_count__i31 (.D(n100[31]), .SP(n7991), .CD(n30648), 
            .CK(debug_c_c), .Q(\register[2][31] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i31.GSR = "ENABLED";
    FD1P3IX uptime_count__i30 (.D(n100[30]), .SP(n7991), .CD(n30648), 
            .CK(debug_c_c), .Q(\register[2][30] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i30.GSR = "ENABLED";
    FD1P3IX uptime_count__i29 (.D(n100[29]), .SP(n7991), .CD(n30649), 
            .CK(debug_c_c), .Q(\register[2][29] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i29.GSR = "ENABLED";
    FD1P3IX uptime_count__i28 (.D(n100[28]), .SP(n7991), .CD(n30649), 
            .CK(debug_c_c), .Q(\register[2][28] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i28.GSR = "ENABLED";
    FD1P3IX uptime_count__i27 (.D(n100[27]), .SP(n7991), .CD(n30649), 
            .CK(debug_c_c), .Q(\register[2][27] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i27.GSR = "ENABLED";
    FD1P3IX uptime_count__i26 (.D(n100[26]), .SP(n7991), .CD(n30649), 
            .CK(debug_c_c), .Q(\register[2][26] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i26.GSR = "ENABLED";
    FD1P3IX uptime_count__i25 (.D(n100[25]), .SP(n7991), .CD(n30649), 
            .CK(debug_c_c), .Q(\register[2][25] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i25.GSR = "ENABLED";
    FD1P3IX uptime_count__i24 (.D(n100[24]), .SP(n7991), .CD(n30649), 
            .CK(debug_c_c), .Q(\register[2][24] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i24.GSR = "ENABLED";
    FD1P3IX uptime_count__i23 (.D(n100[23]), .SP(n7991), .CD(n30649), 
            .CK(debug_c_c), .Q(\register[2][23] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i23.GSR = "ENABLED";
    FD1P3IX uptime_count__i22 (.D(n100[22]), .SP(n7991), .CD(n30648), 
            .CK(debug_c_c), .Q(\register[2][22] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i22.GSR = "ENABLED";
    FD1P3IX uptime_count__i21 (.D(n100[21]), .SP(n7991), .CD(n30648), 
            .CK(debug_c_c), .Q(\register[2][21] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i21.GSR = "ENABLED";
    FD1P3IX uptime_count__i20 (.D(n100[20]), .SP(n7991), .CD(n30648), 
            .CK(debug_c_c), .Q(\register[2][20] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i20.GSR = "ENABLED";
    FD1P3IX uptime_count__i19 (.D(n100[19]), .SP(n7991), .CD(n30648), 
            .CK(debug_c_c), .Q(\register[2][19] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i19.GSR = "ENABLED";
    FD1P3IX uptime_count__i18 (.D(n100[18]), .SP(n7991), .CD(n30648), 
            .CK(debug_c_c), .Q(\register[2][18] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i18.GSR = "ENABLED";
    FD1P3IX uptime_count__i17 (.D(n100[17]), .SP(n7991), .CD(n30648), 
            .CK(debug_c_c), .Q(\register[2][17] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i17.GSR = "ENABLED";
    FD1P3IX uptime_count__i16 (.D(n100[16]), .SP(n7991), .CD(n30648), 
            .CK(debug_c_c), .Q(\register[2][16] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i16.GSR = "ENABLED";
    FD1P3IX uptime_count__i15 (.D(n100[15]), .SP(n7991), .CD(n30648), 
            .CK(debug_c_c), .Q(\register[2][15] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i15.GSR = "ENABLED";
    FD1P3IX uptime_count__i14 (.D(n100[14]), .SP(n7991), .CD(n30649), 
            .CK(debug_c_c), .Q(\register[2][14] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i14.GSR = "ENABLED";
    FD1P3IX uptime_count__i13 (.D(n100[13]), .SP(n7991), .CD(n30648), 
            .CK(debug_c_c), .Q(\register[2][13] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i13.GSR = "ENABLED";
    FD1P3IX uptime_count__i12 (.D(n100[12]), .SP(n7991), .CD(n30649), 
            .CK(debug_c_c), .Q(\register[2][12] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i12.GSR = "ENABLED";
    FD1P3IX uptime_count__i11 (.D(n100[11]), .SP(n7991), .CD(n30649), 
            .CK(debug_c_c), .Q(\register[2][11] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i11.GSR = "ENABLED";
    FD1P3IX uptime_count__i10 (.D(n100[10]), .SP(n7991), .CD(n30649), 
            .CK(debug_c_c), .Q(\register[2][10] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i10.GSR = "ENABLED";
    FD1P3IX uptime_count__i9 (.D(n100[9]), .SP(n7991), .CD(n30649), .CK(debug_c_c), 
            .Q(\register[2][9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i9.GSR = "ENABLED";
    FD1P3IX uptime_count__i8 (.D(n100[8]), .SP(n7991), .CD(n30648), .CK(debug_c_c), 
            .Q(\register[2][8] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i8.GSR = "ENABLED";
    FD1P3IX uptime_count__i7 (.D(n100[7]), .SP(n7991), .CD(n30649), .CK(debug_c_c), 
            .Q(\register[2][7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i7.GSR = "ENABLED";
    FD1P3IX uptime_count__i6 (.D(n100[6]), .SP(n7991), .CD(n30649), .CK(debug_c_c), 
            .Q(\register[2][6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i6.GSR = "ENABLED";
    FD1P3IX uptime_count__i5 (.D(n100[5]), .SP(n7991), .CD(n30648), .CK(debug_c_c), 
            .Q(\register[2][5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i5.GSR = "ENABLED";
    FD1P3IX uptime_count__i4 (.D(n100[4]), .SP(n7991), .CD(n30648), .CK(debug_c_c), 
            .Q(\register[2][4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i4.GSR = "ENABLED";
    FD1P3IX uptime_count__i3 (.D(n100[3]), .SP(n7991), .CD(n30648), .CK(debug_c_c), 
            .Q(\register[2] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i3.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(\register_addr[0] ), .B(n30647), .C(n27213), .D(\select[1] ), 
         .Z(n25733)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut.init = 16'hcdcc;
    FD1P3IX uptime_count__i2 (.D(n100[2]), .SP(n7991), .CD(n28991), .CK(debug_c_c), 
            .Q(\register[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i2.GSR = "ENABLED";
    FD1P3IX uptime_count__i1 (.D(n100[1]), .SP(n7991), .CD(n28991), .CK(debug_c_c), 
            .Q(\register[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i1.GSR = "ENABLED";
    LUT4 i2248_3_lut (.A(prev_clk_1Hz), .B(n30647), .C(clk_1Hz), .Z(n7991)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;
    defparam i2248_3_lut.init = 16'hdcdc;
    LUT4 i114_1_lut (.A(xbee_pause_c), .Z(n178)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(54[26:39])
    defparam i114_1_lut.init = 16'h5555;
    LUT4 i21272_2_lut_rep_262_3_lut_4_lut (.A(\register_addr[5] ), .B(n28972), 
         .C(\register_addr[1] ), .D(\register_addr[2] ), .Z(n28920)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i21272_2_lut_rep_262_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\register_addr[5] ), .B(n28972), .C(n22447), 
         .D(\register_addr[2] ), .Z(n15)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    CCU2D add_134_33 (.A0(\register[2][31] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24232), .S0(n100[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_33.INIT0 = 16'h5aaa;
    defparam add_134_33.INIT1 = 16'h0000;
    defparam add_134_33.INJECT1_0 = "NO";
    defparam add_134_33.INJECT1_1 = "NO";
    CCU2D add_134_31 (.A0(\register[2][29] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][30] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24231), .COUT(n24232), .S0(n100[29]), 
          .S1(n100[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_31.INIT0 = 16'h5aaa;
    defparam add_134_31.INIT1 = 16'h5aaa;
    defparam add_134_31.INJECT1_0 = "NO";
    defparam add_134_31.INJECT1_1 = "NO";
    CCU2D add_134_29 (.A0(\register[2][27] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][28] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24230), .COUT(n24231), .S0(n100[27]), 
          .S1(n100[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_29.INIT0 = 16'h5aaa;
    defparam add_134_29.INIT1 = 16'h5aaa;
    defparam add_134_29.INJECT1_0 = "NO";
    defparam add_134_29.INJECT1_1 = "NO";
    CCU2D add_134_27 (.A0(\register[2][25] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][26] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24229), .COUT(n24230), .S0(n100[25]), 
          .S1(n100[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_27.INIT0 = 16'h5aaa;
    defparam add_134_27.INIT1 = 16'h5aaa;
    defparam add_134_27.INJECT1_0 = "NO";
    defparam add_134_27.INJECT1_1 = "NO";
    CCU2D add_134_25 (.A0(\register[2][23] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][24] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24228), .COUT(n24229), .S0(n100[23]), 
          .S1(n100[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_25.INIT0 = 16'h5aaa;
    defparam add_134_25.INIT1 = 16'h5aaa;
    defparam add_134_25.INJECT1_0 = "NO";
    defparam add_134_25.INJECT1_1 = "NO";
    LUT4 i2_3_lut_3_lut_4_lut (.A(\register_addr[1] ), .B(n28921), .C(n29063), 
         .D(n30647), .Z(n8044)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i2_3_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i20848_2_lut_3_lut_4_lut (.A(\register_addr[1] ), .B(n28921), .C(prev_select), 
         .D(rw), .Z(n27213)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20848_2_lut_3_lut_4_lut.init = 16'hfffe;
    CCU2D add_134_23 (.A0(\register[2][21] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][22] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24227), .COUT(n24228), .S0(n100[21]), 
          .S1(n100[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_23.INIT0 = 16'h5aaa;
    defparam add_134_23.INIT1 = 16'h5aaa;
    defparam add_134_23.INJECT1_0 = "NO";
    defparam add_134_23.INJECT1_1 = "NO";
    CCU2D add_134_21 (.A0(\register[2][19] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][20] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24226), .COUT(n24227), .S0(n100[19]), 
          .S1(n100[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_21.INIT0 = 16'h5aaa;
    defparam add_134_21.INIT1 = 16'h5aaa;
    defparam add_134_21.INJECT1_0 = "NO";
    defparam add_134_21.INJECT1_1 = "NO";
    CCU2D add_134_19 (.A0(\register[2][17] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][18] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24225), .COUT(n24226), .S0(n100[17]), 
          .S1(n100[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_19.INIT0 = 16'h5aaa;
    defparam add_134_19.INIT1 = 16'h5aaa;
    defparam add_134_19.INJECT1_0 = "NO";
    defparam add_134_19.INJECT1_1 = "NO";
    CCU2D add_134_17 (.A0(\register[2][15] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][16] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24224), .COUT(n24225), .S0(n100[15]), 
          .S1(n100[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_17.INIT0 = 16'h5aaa;
    defparam add_134_17.INIT1 = 16'h5aaa;
    defparam add_134_17.INJECT1_0 = "NO";
    defparam add_134_17.INJECT1_1 = "NO";
    CCU2D add_134_15 (.A0(\register[2][13] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][14] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24223), .COUT(n24224), .S0(n100[13]), 
          .S1(n100[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_15.INIT0 = 16'h5aaa;
    defparam add_134_15.INIT1 = 16'h5aaa;
    defparam add_134_15.INJECT1_0 = "NO";
    defparam add_134_15.INJECT1_1 = "NO";
    LUT4 n28059_bdd_2_lut_3_lut_4_lut (.A(n28058), .B(\register_addr[2] ), 
         .C(n29025), .D(n29011), .Z(n28060)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam n28059_bdd_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 n28052_bdd_2_lut_3_lut_4_lut (.A(n28051), .B(\register_addr[2] ), 
         .C(n29025), .D(n29011), .Z(n28053)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam n28052_bdd_2_lut_3_lut_4_lut.init = 16'h0002;
    CCU2D add_134_13 (.A0(\register[2][11] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][12] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24222), .COUT(n24223), .S0(n100[11]), 
          .S1(n100[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_13.INIT0 = 16'h5aaa;
    defparam add_134_13.INIT1 = 16'h5aaa;
    defparam add_134_13.INJECT1_0 = "NO";
    defparam add_134_13.INJECT1_1 = "NO";
    LUT4 register_addr_0__bdd_4_lut_21730 (.A(\register_addr[0] ), .B(\register[2] [1]), 
         .C(\register_addr[1] ), .D(force_pause), .Z(n28051)) /* synthesis lut_function=(!(A (C)+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam register_addr_0__bdd_4_lut_21730.init = 16'h4f4a;
    CCU2D add_134_11 (.A0(\register[2][9] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][10] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24221), .COUT(n24222), .S0(n100[9]), .S1(n100[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_11.INIT0 = 16'h5aaa;
    defparam add_134_11.INIT1 = 16'h5aaa;
    defparam add_134_11.INJECT1_0 = "NO";
    defparam add_134_11.INJECT1_1 = "NO";
    CCU2D add_134_9 (.A0(\register[2][7] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][8] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24220), .COUT(n24221), .S0(n100[7]), .S1(n100[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_9.INIT0 = 16'h5aaa;
    defparam add_134_9.INIT1 = 16'h5aaa;
    defparam add_134_9.INJECT1_0 = "NO";
    defparam add_134_9.INJECT1_1 = "NO";
    CCU2D add_134_7 (.A0(\register[2][5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24219), .COUT(n24220), .S0(n100[5]), .S1(n100[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_7.INIT0 = 16'h5aaa;
    defparam add_134_7.INIT1 = 16'h5aaa;
    defparam add_134_7.INJECT1_0 = "NO";
    defparam add_134_7.INJECT1_1 = "NO";
    CCU2D add_134_5 (.A0(\register[2] [3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2][4] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24218), .COUT(n24219), .S0(n100[3]), .S1(n100[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_5.INIT0 = 16'h5aaa;
    defparam add_134_5.INIT1 = 16'h5aaa;
    defparam add_134_5.INJECT1_0 = "NO";
    defparam add_134_5.INJECT1_1 = "NO";
    CCU2D add_134_3 (.A0(\register[2] [1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24217), .COUT(n24218), .S0(n100[1]), .S1(n100[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_3.INIT0 = 16'h5aaa;
    defparam add_134_3.INIT1 = 16'h5aaa;
    defparam add_134_3.INJECT1_0 = "NO";
    defparam add_134_3.INJECT1_1 = "NO";
    LUT4 \register_0[[2__bdd_4_lut_21719  (.A(\register[0] [2]), .B(\register_addr[1] ), 
         .C(\register[2] [2]), .D(\register_addr[0] ), .Z(n28058)) /* synthesis lut_function=(!(A (B ((D)+!C))+!A (B ((D)+!C)+!B !(D)))) */ ;
    defparam \register_0[[2__bdd_4_lut_21719 .init = 16'h33e2;
    CCU2D add_134_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\register[2] [0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24217), .S1(n100[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_1.INIT0 = 16'hF000;
    defparam add_134_1.INIT1 = 16'h5555;
    defparam add_134_1.INJECT1_0 = "NO";
    defparam add_134_1.INJECT1_1 = "NO";
    LUT4 i885_3_lut (.A(prev_select), .B(n30647), .C(\select[1] ), .Z(n12042)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(61[5] 104[8])
    defparam i885_3_lut.init = 16'h1010;
    LUT4 i21382_2_lut_rep_243_3_lut_4_lut (.A(\register_addr[5] ), .B(n28972), 
         .C(\register_addr[1] ), .D(\register_addr[2] ), .Z(n28901)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i21382_2_lut_rep_243_3_lut_4_lut.init = 16'h0010;
    FD1P3IX read_value__i3 (.D(n6443[3]), .SP(n12042), .CD(n8040), .CK(debug_c_c), 
            .Q(\read_value[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3AX read_value__i4 (.D(n27030), .SP(n12042), .CK(debug_c_c), .Q(\read_value[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3AX read_value__i5 (.D(n27034), .SP(n12042), .CK(debug_c_c), .Q(\read_value[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i5.GSR = "ENABLED";
    LUT4 i14088_4_lut (.A(\register[2] [3]), .B(n48), .C(n11839), .D(n22447), 
         .Z(n6443[3])) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B+(D)))) */ ;
    defparam i14088_4_lut.init = 16'h0a3b;
    FD1P3AX read_value__i6 (.D(n27036), .SP(n12042), .CK(debug_c_c), .Q(\read_value[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i6.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(\register_addr[1] ), .B(n29025), .C(\register_addr[0] ), 
         .D(n28990), .Z(n11839)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i2_4_lut.init = 16'hfffd;
    FD1P3AX read_value__i7 (.D(n27028), .SP(n12042), .CK(debug_c_c), .Q(\read_value[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n27046), .SP(n12042), .CK(debug_c_c), .Q(\read_value[8] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n27042), .SP(n12042), .CK(debug_c_c), .Q(\read_value[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n27045), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[10] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n27026), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[11] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n27025), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[12] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n27027), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[13] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n27029), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[14] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n27038), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[15] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n27031), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[16] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n27033), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[17] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n27023), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[18] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n27041), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[19] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n27047), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[20] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n27048), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[21] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n27040), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[22] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n27039), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[23] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n27035), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[24] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n27050), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[25] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n27024), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[26] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n27049), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[27] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n27044), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[28] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n27032), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[29] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n27037), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[30] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n27043), .SP(n12042), .CK(debug_c_c), 
            .Q(\read_value[31] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n25965), .SP(n12042), .CD(n8040), .CK(debug_c_c), 
            .Q(\read_value[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i0.GSR = "ENABLED";
    FD1P3IX read_size_i0_i1 (.D(n27065), .SP(n12042), .CD(n14380), .CK(debug_c_c), 
            .Q(read_size[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i1.GSR = "ENABLED";
    FD1P3IX read_size_i0_i2 (.D(n15), .SP(n12042), .CD(n14379), .CK(debug_c_c), 
            .Q(read_size[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i2.GSR = "ENABLED";
    FD1P3IX force_pause_151 (.D(\databus[1] ), .SP(n25733), .CD(n28991), 
            .CK(debug_c_c), .Q(force_pause));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam force_pause_151.GSR = "ENABLED";
    LUT4 i3_4_lut (.A(\register_addr[0] ), .B(n28972), .C(\register_addr[5] ), 
         .D(n21_adj_267), .Z(n25965)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i3_4_lut.init = 16'h0100;
    LUT4 i30_4_lut (.A(n29036), .B(\register_addr[1] ), .C(\register_addr[2] ), 
         .D(\register[2] [0]), .Z(n21_adj_267)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam i30_4_lut.init = 16'h3e32;
    \ClockDividerP(factor=12000000)  uptime_div (.GND_net(GND_net), .n30647(n30647), 
            .debug_c_c(debug_c_c), .clk_1Hz(clk_1Hz), .n28991(n28991)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(107[28] 109[53])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000000) 
//

module \ClockDividerP(factor=12000000)  (GND_net, n30647, debug_c_c, clk_1Hz, 
            n28991) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input n30647;
    input debug_c_c;
    output clk_1Hz;
    input n28991;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n24507;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n134;
    
    wire n24506, n24505, n24504, n24503, n24502, n24501, n24500, 
        n24499, n24498, n24497, n24496, n24495, n24494, n24493, 
        n24492, n27500, n2591, n27, n24700, n25, n26, n24, n19, 
        n32, n28, n20, n29, n26_adj_259, n6774, n24601, n24600, 
        n24599, n24598, n24597, n24596, n24595, n24594, n24593, 
        n24592, n24591, n24590;
    
    CCU2D count_2167_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24507), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_33.INIT1 = 16'h0000;
    defparam count_2167_add_4_33.INJECT1_0 = "NO";
    defparam count_2167_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24506), .COUT(n24507), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2167_add_4_31.INJECT1_0 = "NO";
    defparam count_2167_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24505), .COUT(n24506), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2167_add_4_29.INJECT1_0 = "NO";
    defparam count_2167_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24504), .COUT(n24505), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2167_add_4_27.INJECT1_0 = "NO";
    defparam count_2167_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24503), .COUT(n24504), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2167_add_4_25.INJECT1_0 = "NO";
    defparam count_2167_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24502), .COUT(n24503), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2167_add_4_23.INJECT1_0 = "NO";
    defparam count_2167_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24501), .COUT(n24502), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2167_add_4_21.INJECT1_0 = "NO";
    defparam count_2167_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24500), .COUT(n24501), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2167_add_4_19.INJECT1_0 = "NO";
    defparam count_2167_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24499), .COUT(n24500), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2167_add_4_17.INJECT1_0 = "NO";
    defparam count_2167_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24498), .COUT(n24499), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2167_add_4_15.INJECT1_0 = "NO";
    defparam count_2167_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24497), .COUT(n24498), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2167_add_4_13.INJECT1_0 = "NO";
    defparam count_2167_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24496), .COUT(n24497), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2167_add_4_11.INJECT1_0 = "NO";
    defparam count_2167_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24495), .COUT(n24496), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2167_add_4_9.INJECT1_0 = "NO";
    defparam count_2167_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24494), .COUT(n24495), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2167_add_4_7.INJECT1_0 = "NO";
    defparam count_2167_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24493), .COUT(n24494), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2167_add_4_5.INJECT1_0 = "NO";
    defparam count_2167_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24492), .COUT(n24493), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2167_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2167_add_4_3.INJECT1_0 = "NO";
    defparam count_2167_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2167_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24492), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167_add_4_1.INIT0 = 16'hF000;
    defparam count_2167_add_4_1.INIT1 = 16'h0555;
    defparam count_2167_add_4_1.INJECT1_0 = "NO";
    defparam count_2167_add_4_1.INJECT1_1 = "NO";
    LUT4 i21219_2_lut (.A(n27500), .B(n30647), .Z(n2591)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21219_2_lut.init = 16'heeee;
    LUT4 i21217_4_lut (.A(n27), .B(n24700), .C(n25), .D(n26), .Z(n27500)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i21217_4_lut.init = 16'h0004;
    LUT4 i12_4_lut (.A(count[19]), .B(n24), .C(count[8]), .D(count[14]), 
         .Z(n27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(n19), .B(n32), .C(n28), .D(n20), .Z(n24700)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16_4_lut.init = 16'h8000;
    LUT4 i10_4_lut (.A(count[30]), .B(count[22]), .C(count[13]), .D(count[25]), 
         .Z(n25)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i11_4_lut (.A(count[28]), .B(count[15]), .C(count[31]), .D(count[29]), 
         .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut (.A(count[26]), .B(count[24]), .C(count[10]), .D(count[27]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[18]), .B(count[1]), .Z(n19)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i15_4_lut (.A(n29), .B(count[9]), .C(n26_adj_259), .D(count[0]), 
         .Z(n32)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i15_4_lut.init = 16'h8000;
    LUT4 i11_4_lut_adj_258 (.A(count[3]), .B(count[12]), .C(count[5]), 
         .D(count[17]), .Z(n28)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i11_4_lut_adj_258.init = 16'h8000;
    LUT4 i3_2_lut (.A(count[2]), .B(count[11]), .Z(n20)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_259 (.A(count[20]), .B(count[7]), .C(count[23]), 
         .D(count[21]), .Z(n29)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12_4_lut_adj_259.init = 16'h8000;
    LUT4 i9_3_lut (.A(count[16]), .B(count[4]), .C(count[6]), .Z(n26_adj_259)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i9_3_lut.init = 16'h8080;
    FD1S3IX count_2167__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2591), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i0.GSR = "ENABLED";
    FD1S3IX clk_o_14 (.D(n6774), .CK(debug_c_c), .CD(n28991), .Q(clk_1Hz));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D add_18238_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24601), 
          .S0(n6774));
    defparam add_18238_cout.INIT0 = 16'h0000;
    defparam add_18238_cout.INIT1 = 16'h0000;
    defparam add_18238_cout.INJECT1_0 = "NO";
    defparam add_18238_cout.INJECT1_1 = "NO";
    CCU2D add_18238_24 (.A0(count[30]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[31]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24600), .COUT(n24601));
    defparam add_18238_24.INIT0 = 16'h5555;
    defparam add_18238_24.INIT1 = 16'h5555;
    defparam add_18238_24.INJECT1_0 = "NO";
    defparam add_18238_24.INJECT1_1 = "NO";
    CCU2D add_18238_22 (.A0(count[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[29]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24599), .COUT(n24600));
    defparam add_18238_22.INIT0 = 16'h5555;
    defparam add_18238_22.INIT1 = 16'h5555;
    defparam add_18238_22.INJECT1_0 = "NO";
    defparam add_18238_22.INJECT1_1 = "NO";
    CCU2D add_18238_20 (.A0(count[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24598), .COUT(n24599));
    defparam add_18238_20.INIT0 = 16'h5555;
    defparam add_18238_20.INIT1 = 16'h5555;
    defparam add_18238_20.INJECT1_0 = "NO";
    defparam add_18238_20.INJECT1_1 = "NO";
    CCU2D add_18238_18 (.A0(count[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24597), .COUT(n24598));
    defparam add_18238_18.INIT0 = 16'h5555;
    defparam add_18238_18.INIT1 = 16'h5555;
    defparam add_18238_18.INJECT1_0 = "NO";
    defparam add_18238_18.INJECT1_1 = "NO";
    CCU2D add_18238_16 (.A0(count[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24596), .COUT(n24597));
    defparam add_18238_16.INIT0 = 16'h5aaa;
    defparam add_18238_16.INIT1 = 16'h5555;
    defparam add_18238_16.INJECT1_0 = "NO";
    defparam add_18238_16.INJECT1_1 = "NO";
    CCU2D add_18238_14 (.A0(count[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24595), .COUT(n24596));
    defparam add_18238_14.INIT0 = 16'h5aaa;
    defparam add_18238_14.INIT1 = 16'h5555;
    defparam add_18238_14.INJECT1_0 = "NO";
    defparam add_18238_14.INJECT1_1 = "NO";
    CCU2D add_18238_12 (.A0(count[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24594), .COUT(n24595));
    defparam add_18238_12.INIT0 = 16'h5555;
    defparam add_18238_12.INIT1 = 16'h5aaa;
    defparam add_18238_12.INJECT1_0 = "NO";
    defparam add_18238_12.INJECT1_1 = "NO";
    CCU2D add_18238_10 (.A0(count[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24593), .COUT(n24594));
    defparam add_18238_10.INIT0 = 16'h5aaa;
    defparam add_18238_10.INIT1 = 16'h5aaa;
    defparam add_18238_10.INJECT1_0 = "NO";
    defparam add_18238_10.INJECT1_1 = "NO";
    CCU2D add_18238_8 (.A0(count[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24592), .COUT(n24593));
    defparam add_18238_8.INIT0 = 16'h5555;
    defparam add_18238_8.INIT1 = 16'h5aaa;
    defparam add_18238_8.INJECT1_0 = "NO";
    defparam add_18238_8.INJECT1_1 = "NO";
    CCU2D add_18238_6 (.A0(count[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24591), .COUT(n24592));
    defparam add_18238_6.INIT0 = 16'h5555;
    defparam add_18238_6.INIT1 = 16'h5555;
    defparam add_18238_6.INJECT1_0 = "NO";
    defparam add_18238_6.INJECT1_1 = "NO";
    CCU2D add_18238_4 (.A0(count[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24590), .COUT(n24591));
    defparam add_18238_4.INIT0 = 16'h5aaa;
    defparam add_18238_4.INIT1 = 16'h5aaa;
    defparam add_18238_4.INJECT1_0 = "NO";
    defparam add_18238_4.INJECT1_1 = "NO";
    CCU2D add_18238_2 (.A0(count[8]), .B0(count[7]), .C0(GND_net), .D0(GND_net), 
          .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24590));
    defparam add_18238_2.INIT0 = 16'h7000;
    defparam add_18238_2.INIT1 = 16'h5555;
    defparam add_18238_2.INJECT1_0 = "NO";
    defparam add_18238_2.INJECT1_1 = "NO";
    FD1S3IX count_2167__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2591), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i1.GSR = "ENABLED";
    FD1S3IX count_2167__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2591), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i2.GSR = "ENABLED";
    FD1S3IX count_2167__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2591), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i3.GSR = "ENABLED";
    FD1S3IX count_2167__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2591), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i4.GSR = "ENABLED";
    FD1S3IX count_2167__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2591), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i5.GSR = "ENABLED";
    FD1S3IX count_2167__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2591), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i6.GSR = "ENABLED";
    FD1S3IX count_2167__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2591), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i7.GSR = "ENABLED";
    FD1S3IX count_2167__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2591), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i8.GSR = "ENABLED";
    FD1S3IX count_2167__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2591), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i9.GSR = "ENABLED";
    FD1S3IX count_2167__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i10.GSR = "ENABLED";
    FD1S3IX count_2167__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i11.GSR = "ENABLED";
    FD1S3IX count_2167__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i12.GSR = "ENABLED";
    FD1S3IX count_2167__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i13.GSR = "ENABLED";
    FD1S3IX count_2167__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i14.GSR = "ENABLED";
    FD1S3IX count_2167__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i15.GSR = "ENABLED";
    FD1S3IX count_2167__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i16.GSR = "ENABLED";
    FD1S3IX count_2167__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i17.GSR = "ENABLED";
    FD1S3IX count_2167__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i18.GSR = "ENABLED";
    FD1S3IX count_2167__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i19.GSR = "ENABLED";
    FD1S3IX count_2167__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i20.GSR = "ENABLED";
    FD1S3IX count_2167__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i21.GSR = "ENABLED";
    FD1S3IX count_2167__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i22.GSR = "ENABLED";
    FD1S3IX count_2167__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i23.GSR = "ENABLED";
    FD1S3IX count_2167__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i24.GSR = "ENABLED";
    FD1S3IX count_2167__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i25.GSR = "ENABLED";
    FD1S3IX count_2167__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i26.GSR = "ENABLED";
    FD1S3IX count_2167__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i27.GSR = "ENABLED";
    FD1S3IX count_2167__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i28.GSR = "ENABLED";
    FD1S3IX count_2167__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i29.GSR = "ENABLED";
    FD1S3IX count_2167__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i30.GSR = "ENABLED";
    FD1S3IX count_2167__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2591), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2167__i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0110000) 
//

module \ArmPeripheral(axis_haddr=8'b0110000)  (databus, n3176, \register_addr[1] , 
            steps_reg, debug_c_c, n30650, n15, \register_addr[0] , 
            VCC_net, GND_net, Stepper_A_nFault_c, \read_size[0] , n12590, 
            n26777, n14, Stepper_A_M0_c_0, n580, \div_factor_reg[0] , 
            n12230, prev_select, n28946, n28910, n30648, n30649, 
            \div_factor_reg[4] , n609, n611, \control_reg[7] , Stepper_A_Dir_c, 
            \control_reg[4] , Stepper_A_M2_c_2, Stepper_A_M1_c_1, \read_size[2] , 
            n26870, read_value, n28929, n6120, n30651, n30652, \steps_reg[16] , 
            \steps_reg[8] , \steps_reg[5] , \steps_reg[4] , \steps_reg[3] , 
            n26918, stepping, n30647, \div_factor_reg[8] , \div_factor_reg[16] , 
            n17, n7, \select[4] , \register_addr[5] , limit_c_3, Stepper_A_En_c, 
            Stepper_A_Step_c, n24911, n26917, n27444, \register_addr[4] , 
            n11636, n28991) /* synthesis syn_module_defined=1 */ ;
    input [31:0]databus;
    input n3176;
    input \register_addr[1] ;
    output [31:0]steps_reg;
    input debug_c_c;
    input n30650;
    input n15;
    input \register_addr[0] ;
    input VCC_net;
    input GND_net;
    input Stepper_A_nFault_c;
    output \read_size[0] ;
    input n12590;
    input n26777;
    input n14;
    output Stepper_A_M0_c_0;
    input n580;
    output \div_factor_reg[0] ;
    input n12230;
    output prev_select;
    input n28946;
    input n28910;
    input n30648;
    input n30649;
    output \div_factor_reg[4] ;
    input n609;
    input n611;
    output \control_reg[7] ;
    output Stepper_A_Dir_c;
    output \control_reg[4] ;
    output Stepper_A_M2_c_2;
    output Stepper_A_M1_c_1;
    output \read_size[2] ;
    input n26870;
    output [31:0]read_value;
    input n28929;
    input n6120;
    input n30651;
    input n30652;
    output \steps_reg[16] ;
    output \steps_reg[8] ;
    output \steps_reg[5] ;
    output \steps_reg[4] ;
    output \steps_reg[3] ;
    input n26918;
    input stepping;
    input n30647;
    output \div_factor_reg[8] ;
    output \div_factor_reg[16] ;
    input n17;
    input n7;
    input \select[4] ;
    input \register_addr[5] ;
    input limit_c_3;
    output Stepper_A_En_c;
    output Stepper_A_Step_c;
    output n24911;
    input n26917;
    input n27444;
    input \register_addr[4] ;
    output n11636;
    input n28991;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]n225;
    wire [31:0]n3177;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n18790;
    wire [7:0]n7339;
    
    wire n5, n6;
    wire [31:0]n6092;
    
    wire fault_latched, n18787, n18789, n12262, prev_step_clk, step_clk, 
        limit_latched, n183, prev_limit_latched, n12091, n9598;
    wire [31:0]steps_reg_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire int_step, n20613, n28907, n27477, n27474, n26923, n26921, 
        n26925, n26928, n26922, n26920, n26919, n26926, n26927, 
        n26929, n26930, n26931, n26932, n26933, n26934, n26935, 
        n26936, n26937, n26938, n26924, n24372;
    wire [31:0]n6056;
    
    wire n27472, n27473, n24371, n27475, n27476;
    wire [31:0]n100;
    
    wire n24370, n24369, n24368, n24367, n24366, n24365, n24364, 
        n24363, n24362, n24361, n24360, n24359, n24358, n24357, 
        n49, n62_adj_257, n58, n50, n41, n60_adj_258, n54, n42, 
        n52, n38, n56, n46;
    
    LUT4 mux_1310_i1_3_lut (.A(n225[0]), .B(databus[0]), .C(n3176), .Z(n3177[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i1_3_lut.init = 16'hcaca;
    LUT4 i13047_3_lut (.A(control_reg[3]), .B(div_factor_reg[3]), .C(\register_addr[1] ), 
         .Z(n18790)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13047_3_lut.init = 16'hcaca;
    PFUMX i6 (.BLUT(n7339[6]), .ALUT(n5), .C0(\register_addr[1] ), .Z(n6));
    FD1S3IX steps_reg__i0 (.D(n3177[0]), .CK(debug_c_c), .CD(n30650), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    PFUMX i13049 (.BLUT(n18790), .ALUT(n15), .C0(\register_addr[0] ), 
          .Z(n6092[3]));
    IFS1P3DX fault_latched_179 (.D(Stepper_A_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_179.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n26777), .SP(n12590), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    PFUMX i13046 (.BLUT(n18787), .ALUT(n14), .C0(\register_addr[0] ), 
          .Z(n18789));
    FD1P3AX control_reg_i1 (.D(n580), .SP(n12262), .CK(debug_c_c), .Q(Stepper_A_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_176 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_176.GSR = "ENABLED";
    FD1S3AX limit_latched_177 (.D(n183), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_177.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_178 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_178.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n580), .SP(n12230), .CK(debug_c_c), 
            .Q(\div_factor_reg[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_175 (.D(n28946), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_175.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n28910), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n28910), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n28910), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n28910), .PD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n28910), .PD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n28910), .PD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n28910), .PD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n28910), .PD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n28910), .PD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n28910), .PD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n609), .SP(n12230), .CK(debug_c_c), 
            .Q(\div_factor_reg[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n611), .SP(n12230), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n12091), .CD(n9598), .CK(debug_c_c), 
            .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3IX control_reg_i7 (.D(databus[6]), .SP(n12091), .CD(n30649), 
            .CK(debug_c_c), .Q(control_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n12091), .PD(n30649), 
            .CK(debug_c_c), .Q(Stepper_A_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n609), .SP(n12262), .CK(debug_c_c), .Q(\control_reg[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n12091), .PD(n30650), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n611), .SP(n12262), .CK(debug_c_c), .Q(Stepper_A_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n12091), .PD(n30650), 
            .CK(debug_c_c), .Q(Stepper_A_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n26870), .SP(n12590), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3177[31]), .CK(debug_c_c), .CD(n30650), 
            .Q(steps_reg_c[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1P3AX int_step_183 (.D(n28907), .SP(n20613), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_183.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n27477), .SP(n12590), .CD(n28929), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n27474), .SP(n12590), .CD(n28929), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6092[3]), .SP(n12590), .CD(n28929), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6120), .SP(n12590), .CD(n28929), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3177[30]), .CK(debug_c_c), .CD(n30650), 
            .Q(steps_reg_c[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3177[29]), .CK(debug_c_c), .CD(n30650), 
            .Q(steps_reg_c[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3177[28]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg_c[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3177[27]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg_c[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3177[26]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg_c[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3177[25]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg_c[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3177[24]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg_c[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3177[23]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg_c[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3177[22]), .CK(debug_c_c), .CD(n30648), 
            .Q(steps_reg_c[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3177[21]), .CK(debug_c_c), .CD(n30648), 
            .Q(steps_reg_c[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3177[20]), .CK(debug_c_c), .CD(n30648), 
            .Q(steps_reg_c[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3177[19]), .CK(debug_c_c), .CD(n30648), 
            .Q(steps_reg_c[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3177[18]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg_c[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3177[17]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg_c[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3177[16]), .CK(debug_c_c), .CD(n30651), 
            .Q(\steps_reg[16] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3177[15]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg_c[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3177[14]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg_c[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3177[13]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg_c[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3177[12]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg_c[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3177[11]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg_c[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3177[10]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg_c[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3177[9]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg_c[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3177[8]), .CK(debug_c_c), .CD(n30652), 
            .Q(\steps_reg[8] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3177[7]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg_c[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3177[6]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg_c[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3177[5]), .CK(debug_c_c), .CD(n30652), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3177[4]), .CK(debug_c_c), .CD(n30652), 
            .Q(\steps_reg[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3177[3]), .CK(debug_c_c), .CD(n30652), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3177[2]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg_c[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3177[1]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg_c[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n18789), .SP(n12590), .CD(n28929), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6), .SP(n12590), .CD(n28929), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6092[7]), .SP(n12590), .CD(n28929), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n26918), .SP(n12590), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n26923), .SP(n12590), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n26921), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n26925), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n26928), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n26922), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n26920), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n26919), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n26926), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n26927), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n26929), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n26930), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n26931), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n26932), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n26933), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n26934), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    LUT4 i13044_3_lut (.A(Stepper_A_Dir_c), .B(div_factor_reg[5]), .C(\register_addr[1] ), 
         .Z(n18787)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13044_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i27 (.D(n26935), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n26936), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n26937), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n26938), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n26924), .SP(n12590), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    CCU2D sub_126_add_2_33 (.A0(steps_reg_c[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24372), .S0(n225[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_33.INIT0 = 16'h5555;
    defparam sub_126_add_2_33.INIT1 = 16'h0000;
    defparam sub_126_add_2_33.INJECT1_0 = "NO";
    defparam sub_126_add_2_33.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_249 (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .Z(n28907)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i2_3_lut_rep_249.init = 16'h0808;
    LUT4 i14868_4_lut_4_lut (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .D(n30647), .Z(n20613)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i14868_4_lut_4_lut.init = 16'h0038;
    LUT4 i14093_2_lut (.A(\control_reg[7] ), .B(\register_addr[0] ), .Z(n7339[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14093_2_lut.init = 16'h2222;
    LUT4 mux_1668_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg_c[7]), .C(\register_addr[0] ), 
         .Z(n6056[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1668_i8_3_lut.init = 16'hcaca;
    LUT4 i21102_3_lut (.A(Stepper_A_M2_c_2), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n27472)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21102_3_lut.init = 16'hcaca;
    LUT4 i21103_3_lut (.A(div_factor_reg[2]), .B(steps_reg_c[2]), .C(\register_addr[0] ), 
         .Z(n27473)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21103_3_lut.init = 16'hcaca;
    CCU2D sub_126_add_2_31 (.A0(steps_reg_c[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg_c[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24371), .COUT(n24372), .S0(n225[29]), 
          .S1(n225[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_31.INIT0 = 16'h5555;
    defparam sub_126_add_2_31.INIT1 = 16'h5555;
    defparam sub_126_add_2_31.INJECT1_0 = "NO";
    defparam sub_126_add_2_31.INJECT1_1 = "NO";
    LUT4 i21105_3_lut (.A(Stepper_A_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n27475)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21105_3_lut.init = 16'hcaca;
    LUT4 i21106_3_lut (.A(div_factor_reg[1]), .B(steps_reg_c[1]), .C(\register_addr[0] ), 
         .Z(n27476)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21106_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n12230), .CD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n12230), .CD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n12230), .CD(n30649), 
            .CK(debug_c_c), .Q(\div_factor_reg[8] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n12230), .CD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n12230), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n12230), .CD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n12230), .CD(n30649), 
            .CK(debug_c_c), .Q(\div_factor_reg[16] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n12230), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n12230), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n12230), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n12230), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n12230), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n12590), .CD(n28929), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n12590), .CD(n28929), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n17), .SP(n12590), .CD(n28929), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    LUT4 i21310_2_lut (.A(n12091), .B(n30647), .Z(n12262)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21310_2_lut.init = 16'heeee;
    LUT4 i21237_4_lut (.A(n7), .B(\select[4] ), .C(\register_addr[5] ), 
         .D(prev_select), .Z(n12091)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i21237_4_lut.init = 16'h0040;
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n12230), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    CCU2D sub_126_add_2_29 (.A0(steps_reg_c[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg_c[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24370), .COUT(n24371), .S0(n225[27]), 
          .S1(n225[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_29.INIT0 = 16'h5555;
    defparam sub_126_add_2_29.INIT1 = 16'h5555;
    defparam sub_126_add_2_29.INJECT1_0 = "NO";
    defparam sub_126_add_2_29.INJECT1_1 = "NO";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n12230), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n12230), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    LUT4 i119_1_lut (.A(limit_c_3), .Z(n183)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i119_1_lut.init = 16'h5555;
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n12230), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n12230), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n12230), .CD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n12230), .CD(n30649), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    LUT4 i8_1_lut (.A(control_reg[6]), .Z(Stepper_A_En_c)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(44[14:29])
    defparam i8_1_lut.init = 16'h5555;
    LUT4 i21206_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_A_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i21206_2_lut.init = 16'h9999;
    CCU2D sub_126_add_2_27 (.A0(steps_reg_c[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg_c[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24369), .COUT(n24370), .S0(n225[25]), 
          .S1(n225[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_27.INIT0 = 16'h5555;
    defparam sub_126_add_2_27.INIT1 = 16'h5555;
    defparam sub_126_add_2_27.INJECT1_0 = "NO";
    defparam sub_126_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_25 (.A0(steps_reg_c[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg_c[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24368), .COUT(n24369), .S0(n225[23]), 
          .S1(n225[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_25.INIT0 = 16'h5555;
    defparam sub_126_add_2_25.INIT1 = 16'h5555;
    defparam sub_126_add_2_25.INJECT1_0 = "NO";
    defparam sub_126_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_23 (.A0(steps_reg_c[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg_c[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24367), .COUT(n24368), .S0(n225[21]), 
          .S1(n225[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_23.INIT0 = 16'h5555;
    defparam sub_126_add_2_23.INIT1 = 16'h5555;
    defparam sub_126_add_2_23.INJECT1_0 = "NO";
    defparam sub_126_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_21 (.A0(steps_reg_c[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg_c[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24366), .COUT(n24367), .S0(n225[19]), 
          .S1(n225[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_21.INIT0 = 16'h5555;
    defparam sub_126_add_2_21.INIT1 = 16'h5555;
    defparam sub_126_add_2_21.INJECT1_0 = "NO";
    defparam sub_126_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_19 (.A0(steps_reg_c[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg_c[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24365), .COUT(n24366), .S0(n225[17]), 
          .S1(n225[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_19.INIT0 = 16'h5555;
    defparam sub_126_add_2_19.INIT1 = 16'h5555;
    defparam sub_126_add_2_19.INJECT1_0 = "NO";
    defparam sub_126_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_17 (.A0(steps_reg_c[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[16] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24364), .COUT(n24365), .S0(n225[15]), 
          .S1(n225[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_17.INIT0 = 16'h5555;
    defparam sub_126_add_2_17.INIT1 = 16'h5555;
    defparam sub_126_add_2_17.INJECT1_0 = "NO";
    defparam sub_126_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_15 (.A0(steps_reg_c[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg_c[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24363), .COUT(n24364), .S0(n225[13]), 
          .S1(n225[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_15.INIT0 = 16'h5555;
    defparam sub_126_add_2_15.INIT1 = 16'h5555;
    defparam sub_126_add_2_15.INJECT1_0 = "NO";
    defparam sub_126_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_13 (.A0(steps_reg_c[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg_c[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24362), .COUT(n24363), .S0(n225[11]), 
          .S1(n225[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_13.INIT0 = 16'h5555;
    defparam sub_126_add_2_13.INIT1 = 16'h5555;
    defparam sub_126_add_2_13.INJECT1_0 = "NO";
    defparam sub_126_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_11 (.A0(steps_reg_c[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg_c[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24361), .COUT(n24362), .S0(n225[9]), .S1(n225[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_11.INIT0 = 16'h5555;
    defparam sub_126_add_2_11.INIT1 = 16'h5555;
    defparam sub_126_add_2_11.INJECT1_0 = "NO";
    defparam sub_126_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_9 (.A0(steps_reg_c[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[8] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24360), .COUT(n24361), .S0(n225[7]), .S1(n225[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_9.INIT0 = 16'h5555;
    defparam sub_126_add_2_9.INIT1 = 16'h5555;
    defparam sub_126_add_2_9.INJECT1_0 = "NO";
    defparam sub_126_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg_c[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24359), .COUT(n24360), .S0(n225[5]), .S1(n225[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_7.INIT0 = 16'h5555;
    defparam sub_126_add_2_7.INIT1 = 16'h5555;
    defparam sub_126_add_2_7.INJECT1_0 = "NO";
    defparam sub_126_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[4] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24358), .COUT(n24359), .S0(n225[3]), .S1(n225[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_5.INIT0 = 16'h5555;
    defparam sub_126_add_2_5.INIT1 = 16'h5555;
    defparam sub_126_add_2_5.INJECT1_0 = "NO";
    defparam sub_126_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_3 (.A0(steps_reg_c[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg_c[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24357), .COUT(n24358), .S0(n225[1]), .S1(n225[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_3.INIT0 = 16'h5555;
    defparam sub_126_add_2_3.INIT1 = 16'h5555;
    defparam sub_126_add_2_3.INJECT1_0 = "NO";
    defparam sub_126_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(stepping), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n24357), .S1(n225[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_1.INIT0 = 16'h0000;
    defparam sub_126_add_2_1.INIT1 = 16'h5595;
    defparam sub_126_add_2_1.INJECT1_0 = "NO";
    defparam sub_126_add_2_1.INJECT1_1 = "NO";
    LUT4 i3837_3_lut (.A(prev_limit_latched), .B(n30647), .C(limit_latched), 
         .Z(n9598)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i3837_3_lut.init = 16'hdcdc;
    LUT4 mux_1310_i32_3_lut (.A(n225[31]), .B(databus[31]), .C(n3176), 
         .Z(n3177[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i32_3_lut.init = 16'hcaca;
    LUT4 i14094_2_lut (.A(control_reg[6]), .B(\register_addr[0] ), .Z(n7339[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14094_2_lut.init = 16'h2222;
    LUT4 i5_3_lut (.A(div_factor_reg[6]), .B(steps_reg_c[6]), .C(\register_addr[0] ), 
         .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i5_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62_adj_257), .C(n58), .D(n50), .Z(n24911)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[0]), .B(steps_reg_c[9]), .C(steps_reg_c[28]), 
         .D(steps_reg_c[2]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut (.A(div_factor_reg[29]), .B(n26917), .C(steps_reg_c[29]), 
         .D(\register_addr[0] ), .Z(n26937)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i30_4_lut (.A(n41), .B(n60_adj_258), .C(n54), .D(n42), .Z(n62_adj_257)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg_c[25]), .B(n52), .C(n38), .D(steps_reg_c[26]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(\steps_reg[4] ), .B(steps_reg_c[11]), .C(\steps_reg[16] ), 
         .D(steps_reg_c[21]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg_c[30]), .B(steps_reg_c[7]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg_c[20]), .B(n56), .C(n46), .D(steps_reg_c[15]), 
         .Z(n60_adj_258)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg_c[22]), .B(steps_reg_c[12]), .C(steps_reg_c[6]), 
         .D(steps_reg_c[18]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg_c[14]), .B(steps_reg_c[19]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg_c[13]), .B(steps_reg_c[17]), .C(\steps_reg[5] ), 
         .D(steps_reg_c[31]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg_c[23]), .B(steps_reg_c[29]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_239 (.A(div_factor_reg[30]), .B(n26917), .C(steps_reg_c[30]), 
         .D(\register_addr[0] ), .Z(n26938)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_239.init = 16'hc088;
    LUT4 i1_4_lut_adj_240 (.A(div_factor_reg[31]), .B(n26917), .C(steps_reg_c[31]), 
         .D(\register_addr[0] ), .Z(n26924)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_240.init = 16'hc088;
    LUT4 i20_4_lut (.A(steps_reg_c[24]), .B(\steps_reg[8] ), .C(steps_reg_c[1]), 
         .D(steps_reg_c[27]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg_c[10]), .B(\steps_reg[3] ), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 mux_1310_i31_3_lut (.A(n225[30]), .B(databus[30]), .C(n3176), 
         .Z(n3177[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i30_3_lut (.A(n225[29]), .B(databus[29]), .C(n3176), 
         .Z(n3177[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i29_3_lut (.A(n225[28]), .B(databus[28]), .C(n3176), 
         .Z(n3177[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i28_3_lut (.A(n225[27]), .B(databus[27]), .C(n3176), 
         .Z(n3177[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i27_3_lut (.A(n225[26]), .B(databus[26]), .C(n3176), 
         .Z(n3177[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i26_3_lut (.A(n225[25]), .B(databus[25]), .C(n3176), 
         .Z(n3177[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i25_3_lut (.A(n225[24]), .B(databus[24]), .C(n3176), 
         .Z(n3177[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i24_3_lut (.A(n225[23]), .B(databus[23]), .C(n3176), 
         .Z(n3177[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i23_3_lut (.A(n225[22]), .B(databus[22]), .C(n3176), 
         .Z(n3177[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i22_3_lut (.A(n225[21]), .B(databus[21]), .C(n3176), 
         .Z(n3177[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i21_3_lut (.A(n225[20]), .B(databus[20]), .C(n3176), 
         .Z(n3177[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i20_3_lut (.A(n225[19]), .B(databus[19]), .C(n3176), 
         .Z(n3177[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i19_3_lut (.A(n225[18]), .B(databus[18]), .C(n3176), 
         .Z(n3177[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i18_3_lut (.A(n225[17]), .B(databus[17]), .C(n3176), 
         .Z(n3177[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i17_3_lut (.A(n225[16]), .B(databus[16]), .C(n3176), 
         .Z(n3177[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i16_3_lut (.A(n225[15]), .B(databus[15]), .C(n3176), 
         .Z(n3177[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i15_3_lut (.A(n225[14]), .B(databus[14]), .C(n3176), 
         .Z(n3177[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i14_3_lut (.A(n225[13]), .B(databus[13]), .C(n3176), 
         .Z(n3177[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i13_3_lut (.A(n225[12]), .B(databus[12]), .C(n3176), 
         .Z(n3177[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i12_3_lut (.A(n225[11]), .B(databus[11]), .C(n3176), 
         .Z(n3177[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i11_3_lut (.A(n225[10]), .B(databus[10]), .C(n3176), 
         .Z(n3177[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i10_3_lut (.A(n225[9]), .B(databus[9]), .C(n3176), .Z(n3177[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i9_3_lut (.A(n225[8]), .B(databus[8]), .C(n3176), .Z(n3177[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i8_3_lut (.A(n225[7]), .B(databus[7]), .C(n3176), .Z(n3177[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i7_3_lut (.A(n225[6]), .B(databus[6]), .C(n3176), .Z(n3177[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i6_3_lut (.A(n225[5]), .B(databus[5]), .C(n3176), .Z(n3177[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i5_3_lut (.A(n225[4]), .B(databus[4]), .C(n3176), .Z(n3177[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i4_3_lut (.A(n225[3]), .B(databus[3]), .C(n3176), .Z(n3177[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i3_3_lut (.A(n225[2]), .B(databus[2]), .C(n3176), .Z(n3177[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1310_i2_3_lut (.A(n225[1]), .B(databus[1]), .C(n3176), .Z(n3177[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1310_i2_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i0 (.D(n27444), .SP(n12590), .CD(n28929), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    PFUMX mux_1672_i8 (.BLUT(n7339[7]), .ALUT(n6056[7]), .C0(\register_addr[1] ), 
          .Z(n6092[7]));
    PFUMX i21104 (.BLUT(n27472), .ALUT(n27473), .C0(\register_addr[1] ), 
          .Z(n27474));
    PFUMX i21107 (.BLUT(n27475), .ALUT(n27476), .C0(\register_addr[1] ), 
          .Z(n27477));
    LUT4 i1_4_lut_adj_241 (.A(div_factor_reg[9]), .B(n26917), .C(steps_reg_c[9]), 
         .D(\register_addr[0] ), .Z(n26923)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_241.init = 16'hc088;
    LUT4 i1_4_lut_adj_242 (.A(div_factor_reg[10]), .B(n26917), .C(steps_reg_c[10]), 
         .D(\register_addr[0] ), .Z(n26921)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_242.init = 16'hc088;
    LUT4 i1_4_lut_adj_243 (.A(div_factor_reg[11]), .B(n26917), .C(steps_reg_c[11]), 
         .D(\register_addr[0] ), .Z(n26925)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_243.init = 16'hc088;
    LUT4 i1_4_lut_adj_244 (.A(div_factor_reg[12]), .B(n26917), .C(steps_reg_c[12]), 
         .D(\register_addr[0] ), .Z(n26928)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_244.init = 16'hc088;
    LUT4 i1_4_lut_adj_245 (.A(div_factor_reg[13]), .B(n26917), .C(steps_reg_c[13]), 
         .D(\register_addr[0] ), .Z(n26922)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_245.init = 16'hc088;
    LUT4 i1_4_lut_adj_246 (.A(div_factor_reg[14]), .B(n26917), .C(steps_reg_c[14]), 
         .D(\register_addr[0] ), .Z(n26920)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_246.init = 16'hc088;
    LUT4 i1_4_lut_adj_247 (.A(div_factor_reg[15]), .B(n26917), .C(steps_reg_c[15]), 
         .D(\register_addr[0] ), .Z(n26919)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_247.init = 16'hc088;
    LUT4 i14090_4_lut (.A(div_factor_reg[18]), .B(\register_addr[1] ), .C(steps_reg_c[18]), 
         .D(\register_addr[0] ), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14090_4_lut.init = 16'hc088;
    LUT4 i14091_4_lut (.A(div_factor_reg[17]), .B(\register_addr[1] ), .C(steps_reg_c[17]), 
         .D(\register_addr[0] ), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14091_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_248 (.A(div_factor_reg[19]), .B(n26917), .C(steps_reg_c[19]), 
         .D(\register_addr[0] ), .Z(n26926)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_248.init = 16'hc088;
    LUT4 i1_4_lut_adj_249 (.A(div_factor_reg[20]), .B(n26917), .C(steps_reg_c[20]), 
         .D(\register_addr[0] ), .Z(n26927)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_249.init = 16'hc088;
    LUT4 i1_2_lut (.A(\register_addr[4] ), .B(\register_addr[5] ), .Z(n11636)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_250 (.A(div_factor_reg[21]), .B(n26917), .C(steps_reg_c[21]), 
         .D(\register_addr[0] ), .Z(n26929)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_250.init = 16'hc088;
    LUT4 i1_4_lut_adj_251 (.A(div_factor_reg[22]), .B(n26917), .C(steps_reg_c[22]), 
         .D(\register_addr[0] ), .Z(n26930)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_251.init = 16'hc088;
    LUT4 i1_4_lut_adj_252 (.A(div_factor_reg[23]), .B(n26917), .C(steps_reg_c[23]), 
         .D(\register_addr[0] ), .Z(n26931)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_252.init = 16'hc088;
    LUT4 i1_4_lut_adj_253 (.A(div_factor_reg[24]), .B(n26917), .C(steps_reg_c[24]), 
         .D(\register_addr[0] ), .Z(n26932)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_253.init = 16'hc088;
    LUT4 i1_4_lut_adj_254 (.A(div_factor_reg[25]), .B(n26917), .C(steps_reg_c[25]), 
         .D(\register_addr[0] ), .Z(n26933)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_254.init = 16'hc088;
    LUT4 i1_4_lut_adj_255 (.A(div_factor_reg[26]), .B(n26917), .C(steps_reg_c[26]), 
         .D(\register_addr[0] ), .Z(n26934)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_255.init = 16'hc088;
    LUT4 i1_4_lut_adj_256 (.A(div_factor_reg[27]), .B(n26917), .C(steps_reg_c[27]), 
         .D(\register_addr[0] ), .Z(n26935)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_256.init = 16'hc088;
    LUT4 i1_4_lut_adj_257 (.A(div_factor_reg[28]), .B(n26917), .C(steps_reg_c[28]), 
         .D(\register_addr[0] ), .Z(n26936)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_257.init = 16'hc088;
    ClockDivider_U9 step_clk_gen (.GND_net(GND_net), .n30647(n30647), .div_factor_reg({div_factor_reg[31:17], 
            \div_factor_reg[16] , div_factor_reg[15:9], \div_factor_reg[8] , 
            div_factor_reg[7:5], \div_factor_reg[4] , div_factor_reg[3:1], 
            \div_factor_reg[0] }), .step_clk(step_clk), .debug_c_c(debug_c_c), 
            .n28991(n28991)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U9
//

module ClockDivider_U9 (GND_net, n30647, div_factor_reg, step_clk, debug_c_c, 
            n28991) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input n30647;
    input [31:0]div_factor_reg;
    output step_clk;
    input debug_c_c;
    input n28991;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n24259;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n40;
    
    wire n24260, n24258, n24257, n24256, n23962;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n23963, n24255, n23961, n24254, n24253, n7156, n28890, 
        n24248, n7190, n24247, n23975, n23976, n24246, n23974, 
        n24245, n24244, n24243, n24242, n7121, n24241, n24240, 
        n23965, n23966, n23964, n23973, n24239, n24238, n24237, 
        n24236, n23972, n24491;
    wire [31:0]n134;
    
    wire n24490, n24235, n24489, n24488, n24234, n24233, n24487, 
        n24486, n24485, n24484, n14388, n24483, n24482, n24481, 
        n24480, n24479, n24478, n24477, n24476, n23971, n24308, 
        n24307, n24306, n24305, n24304, n24303, n24302, n24301, 
        n24300, n24299, n24298, n24297, n24296, n24295, n24294, 
        n24293, n23970, n23969, n23968, n23967, n24268, n24267, 
        n24266, n24265, n24264, n24263, n24262, n24261;
    
    CCU2D sub_1727_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24259), .COUT(n24260));
    defparam sub_1727_add_2_15.INIT0 = 16'h5999;
    defparam sub_1727_add_2_15.INIT1 = 16'h5999;
    defparam sub_1727_add_2_15.INJECT1_0 = "NO";
    defparam sub_1727_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24258), .COUT(n24259));
    defparam sub_1727_add_2_13.INIT0 = 16'h5999;
    defparam sub_1727_add_2_13.INIT1 = 16'h5999;
    defparam sub_1727_add_2_13.INJECT1_0 = "NO";
    defparam sub_1727_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24257), .COUT(n24258));
    defparam sub_1727_add_2_11.INIT0 = 16'h5999;
    defparam sub_1727_add_2_11.INIT1 = 16'h5999;
    defparam sub_1727_add_2_11.INJECT1_0 = "NO";
    defparam sub_1727_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24256), .COUT(n24257));
    defparam sub_1727_add_2_9.INIT0 = 16'h5999;
    defparam sub_1727_add_2_9.INIT1 = 16'h5999;
    defparam sub_1727_add_2_9.INJECT1_0 = "NO";
    defparam sub_1727_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1725_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23962), .COUT(n23963));
    defparam sub_1725_add_2_5.INIT0 = 16'h5999;
    defparam sub_1725_add_2_5.INIT1 = 16'h5999;
    defparam sub_1725_add_2_5.INJECT1_0 = "NO";
    defparam sub_1725_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24255), .COUT(n24256));
    defparam sub_1727_add_2_7.INIT0 = 16'h5999;
    defparam sub_1727_add_2_7.INIT1 = 16'h5999;
    defparam sub_1727_add_2_7.INJECT1_0 = "NO";
    defparam sub_1727_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1725_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23961), .COUT(n23962));
    defparam sub_1725_add_2_3.INIT0 = 16'h5999;
    defparam sub_1725_add_2_3.INIT1 = 16'h5999;
    defparam sub_1725_add_2_3.INJECT1_0 = "NO";
    defparam sub_1725_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24254), .COUT(n24255));
    defparam sub_1727_add_2_5.INIT0 = 16'h5999;
    defparam sub_1727_add_2_5.INIT1 = 16'h5999;
    defparam sub_1727_add_2_5.INJECT1_0 = "NO";
    defparam sub_1727_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24253), .COUT(n24254));
    defparam sub_1727_add_2_3.INIT0 = 16'h5999;
    defparam sub_1727_add_2_3.INIT1 = 16'h5999;
    defparam sub_1727_add_2_3.INJECT1_0 = "NO";
    defparam sub_1727_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n24253));
    defparam sub_1727_add_2_1.INIT0 = 16'h0000;
    defparam sub_1727_add_2_1.INIT1 = 16'h5999;
    defparam sub_1727_add_2_1.INJECT1_0 = "NO";
    defparam sub_1727_add_2_1.INJECT1_1 = "NO";
    LUT4 i962_2_lut_rep_232 (.A(n7156), .B(n30647), .Z(n28890)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i962_2_lut_rep_232.init = 16'heeee;
    CCU2D sub_1728_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24248), .S1(n7190));
    defparam sub_1728_add_2_33.INIT0 = 16'hf555;
    defparam sub_1728_add_2_33.INIT1 = 16'h0000;
    defparam sub_1728_add_2_33.INJECT1_0 = "NO";
    defparam sub_1728_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1728_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24247), .COUT(n24248));
    defparam sub_1728_add_2_31.INIT0 = 16'hf555;
    defparam sub_1728_add_2_31.INIT1 = 16'hf555;
    defparam sub_1728_add_2_31.INJECT1_0 = "NO";
    defparam sub_1728_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1725_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23975), .COUT(n23976));
    defparam sub_1725_add_2_31.INIT0 = 16'h5999;
    defparam sub_1725_add_2_31.INIT1 = 16'h5999;
    defparam sub_1725_add_2_31.INJECT1_0 = "NO";
    defparam sub_1725_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1728_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24246), .COUT(n24247));
    defparam sub_1728_add_2_29.INIT0 = 16'hf555;
    defparam sub_1728_add_2_29.INIT1 = 16'hf555;
    defparam sub_1728_add_2_29.INJECT1_0 = "NO";
    defparam sub_1728_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1725_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23974), .COUT(n23975));
    defparam sub_1725_add_2_29.INIT0 = 16'h5999;
    defparam sub_1725_add_2_29.INIT1 = 16'h5999;
    defparam sub_1725_add_2_29.INJECT1_0 = "NO";
    defparam sub_1725_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1728_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24245), .COUT(n24246));
    defparam sub_1728_add_2_27.INIT0 = 16'hf555;
    defparam sub_1728_add_2_27.INIT1 = 16'hf555;
    defparam sub_1728_add_2_27.INJECT1_0 = "NO";
    defparam sub_1728_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1728_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24244), .COUT(n24245));
    defparam sub_1728_add_2_25.INIT0 = 16'hf555;
    defparam sub_1728_add_2_25.INIT1 = 16'hf555;
    defparam sub_1728_add_2_25.INJECT1_0 = "NO";
    defparam sub_1728_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1728_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24243), .COUT(n24244));
    defparam sub_1728_add_2_23.INIT0 = 16'hf555;
    defparam sub_1728_add_2_23.INIT1 = 16'hf555;
    defparam sub_1728_add_2_23.INJECT1_0 = "NO";
    defparam sub_1728_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1728_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24242), .COUT(n24243));
    defparam sub_1728_add_2_21.INIT0 = 16'hf555;
    defparam sub_1728_add_2_21.INIT1 = 16'hf555;
    defparam sub_1728_add_2_21.INJECT1_0 = "NO";
    defparam sub_1728_add_2_21.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n7121), .CK(debug_c_c), .CD(n28991), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_1728_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24241), .COUT(n24242));
    defparam sub_1728_add_2_19.INIT0 = 16'hf555;
    defparam sub_1728_add_2_19.INIT1 = 16'hf555;
    defparam sub_1728_add_2_19.INJECT1_0 = "NO";
    defparam sub_1728_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1728_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24240), .COUT(n24241));
    defparam sub_1728_add_2_17.INIT0 = 16'hf555;
    defparam sub_1728_add_2_17.INIT1 = 16'hf555;
    defparam sub_1728_add_2_17.INJECT1_0 = "NO";
    defparam sub_1728_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1725_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23965), .COUT(n23966));
    defparam sub_1725_add_2_11.INIT0 = 16'h5999;
    defparam sub_1725_add_2_11.INIT1 = 16'h5999;
    defparam sub_1725_add_2_11.INJECT1_0 = "NO";
    defparam sub_1725_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1725_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23964), .COUT(n23965));
    defparam sub_1725_add_2_9.INIT0 = 16'h5999;
    defparam sub_1725_add_2_9.INIT1 = 16'h5999;
    defparam sub_1725_add_2_9.INJECT1_0 = "NO";
    defparam sub_1725_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1725_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23973), .COUT(n23974));
    defparam sub_1725_add_2_27.INIT0 = 16'h5999;
    defparam sub_1725_add_2_27.INIT1 = 16'h5999;
    defparam sub_1725_add_2_27.INJECT1_0 = "NO";
    defparam sub_1725_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1728_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24239), .COUT(n24240));
    defparam sub_1728_add_2_15.INIT0 = 16'hf555;
    defparam sub_1728_add_2_15.INIT1 = 16'hf555;
    defparam sub_1728_add_2_15.INJECT1_0 = "NO";
    defparam sub_1728_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1728_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24238), .COUT(n24239));
    defparam sub_1728_add_2_13.INIT0 = 16'hf555;
    defparam sub_1728_add_2_13.INIT1 = 16'hf555;
    defparam sub_1728_add_2_13.INJECT1_0 = "NO";
    defparam sub_1728_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1728_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24237), .COUT(n24238));
    defparam sub_1728_add_2_11.INIT0 = 16'hf555;
    defparam sub_1728_add_2_11.INIT1 = 16'hf555;
    defparam sub_1728_add_2_11.INJECT1_0 = "NO";
    defparam sub_1728_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1728_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24236), .COUT(n24237));
    defparam sub_1728_add_2_9.INIT0 = 16'hf555;
    defparam sub_1728_add_2_9.INIT1 = 16'hf555;
    defparam sub_1728_add_2_9.INJECT1_0 = "NO";
    defparam sub_1728_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1725_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23972), .COUT(n23973));
    defparam sub_1725_add_2_25.INIT0 = 16'h5999;
    defparam sub_1725_add_2_25.INIT1 = 16'h5999;
    defparam sub_1725_add_2_25.INJECT1_0 = "NO";
    defparam sub_1725_add_2_25.INJECT1_1 = "NO";
    CCU2D count_2171_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24491), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_33.INIT1 = 16'h0000;
    defparam count_2171_add_4_33.INJECT1_0 = "NO";
    defparam count_2171_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2171_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24490), .COUT(n24491), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2171_add_4_31.INJECT1_0 = "NO";
    defparam count_2171_add_4_31.INJECT1_1 = "NO";
    CCU2D sub_1728_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24235), .COUT(n24236));
    defparam sub_1728_add_2_7.INIT0 = 16'hf555;
    defparam sub_1728_add_2_7.INIT1 = 16'hf555;
    defparam sub_1728_add_2_7.INJECT1_0 = "NO";
    defparam sub_1728_add_2_7.INJECT1_1 = "NO";
    CCU2D count_2171_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24489), .COUT(n24490), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2171_add_4_29.INJECT1_0 = "NO";
    defparam count_2171_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2171_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24488), .COUT(n24489), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2171_add_4_27.INJECT1_0 = "NO";
    defparam count_2171_add_4_27.INJECT1_1 = "NO";
    CCU2D sub_1728_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24234), .COUT(n24235));
    defparam sub_1728_add_2_5.INIT0 = 16'hf555;
    defparam sub_1728_add_2_5.INIT1 = 16'hf555;
    defparam sub_1728_add_2_5.INJECT1_0 = "NO";
    defparam sub_1728_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1728_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24233), .COUT(n24234));
    defparam sub_1728_add_2_3.INIT0 = 16'hf555;
    defparam sub_1728_add_2_3.INIT1 = 16'hf555;
    defparam sub_1728_add_2_3.INJECT1_0 = "NO";
    defparam sub_1728_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1728_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n24233));
    defparam sub_1728_add_2_1.INIT0 = 16'h0000;
    defparam sub_1728_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1728_add_2_1.INJECT1_0 = "NO";
    defparam sub_1728_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2171_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24487), .COUT(n24488), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2171_add_4_25.INJECT1_0 = "NO";
    defparam count_2171_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2171_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24486), .COUT(n24487), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2171_add_4_23.INJECT1_0 = "NO";
    defparam count_2171_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2171_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24485), .COUT(n24486), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2171_add_4_21.INJECT1_0 = "NO";
    defparam count_2171_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2171_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24484), .COUT(n24485), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2171_add_4_19.INJECT1_0 = "NO";
    defparam count_2171_add_4_19.INJECT1_1 = "NO";
    LUT4 i8622_2_lut_3_lut (.A(n7156), .B(n30647), .C(n7190), .Z(n14388)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i8622_2_lut_3_lut.init = 16'he0e0;
    CCU2D count_2171_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24483), .COUT(n24484), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2171_add_4_17.INJECT1_0 = "NO";
    defparam count_2171_add_4_17.INJECT1_1 = "NO";
    FD1S3IX count_2171__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i0.GSR = "ENABLED";
    CCU2D count_2171_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24482), .COUT(n24483), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2171_add_4_15.INJECT1_0 = "NO";
    defparam count_2171_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2171_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24481), .COUT(n24482), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2171_add_4_13.INJECT1_0 = "NO";
    defparam count_2171_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2171_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24480), .COUT(n24481), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2171_add_4_11.INJECT1_0 = "NO";
    defparam count_2171_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2171_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24479), .COUT(n24480), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2171_add_4_9.INJECT1_0 = "NO";
    defparam count_2171_add_4_9.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    CCU2D count_2171_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24478), .COUT(n24479), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2171_add_4_7.INJECT1_0 = "NO";
    defparam count_2171_add_4_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    CCU2D count_2171_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24477), .COUT(n24478), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2171_add_4_5.INJECT1_0 = "NO";
    defparam count_2171_add_4_5.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    CCU2D count_2171_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24476), .COUT(n24477), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2171_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2171_add_4_3.INJECT1_0 = "NO";
    defparam count_2171_add_4_3.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    CCU2D count_2171_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24476), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171_add_4_1.INIT0 = 16'hF000;
    defparam count_2171_add_4_1.INIT1 = 16'h0555;
    defparam count_2171_add_4_1.INJECT1_0 = "NO";
    defparam count_2171_add_4_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    CCU2D sub_1725_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23971), .COUT(n23972));
    defparam sub_1725_add_2_23.INIT0 = 16'h5999;
    defparam sub_1725_add_2_23.INIT1 = 16'h5999;
    defparam sub_1725_add_2_23.INJECT1_0 = "NO";
    defparam sub_1725_add_2_23.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n28890), .PD(n14388), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24308), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24307), .COUT(n24308), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24306), .COUT(n24307), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24305), .COUT(n24306), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24304), .COUT(n24305), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24303), .COUT(n24304), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    FD1S3IX count_2171__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i1.GSR = "ENABLED";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24302), .COUT(n24303), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24301), .COUT(n24302), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24300), .COUT(n24301), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    FD1S3IX count_2171__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i2.GSR = "ENABLED";
    FD1S3IX count_2171__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i3.GSR = "ENABLED";
    FD1S3IX count_2171__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i4.GSR = "ENABLED";
    FD1S3IX count_2171__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i5.GSR = "ENABLED";
    FD1S3IX count_2171__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i6.GSR = "ENABLED";
    FD1S3IX count_2171__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i7.GSR = "ENABLED";
    FD1S3IX count_2171__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i8.GSR = "ENABLED";
    FD1S3IX count_2171__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i9.GSR = "ENABLED";
    FD1S3IX count_2171__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i10.GSR = "ENABLED";
    FD1S3IX count_2171__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i11.GSR = "ENABLED";
    FD1S3IX count_2171__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i12.GSR = "ENABLED";
    FD1S3IX count_2171__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i13.GSR = "ENABLED";
    FD1S3IX count_2171__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i14.GSR = "ENABLED";
    FD1S3IX count_2171__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i15.GSR = "ENABLED";
    FD1S3IX count_2171__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i16.GSR = "ENABLED";
    FD1S3IX count_2171__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i17.GSR = "ENABLED";
    FD1S3IX count_2171__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i18.GSR = "ENABLED";
    FD1S3IX count_2171__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i19.GSR = "ENABLED";
    FD1S3IX count_2171__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i20.GSR = "ENABLED";
    FD1S3IX count_2171__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i21.GSR = "ENABLED";
    FD1S3IX count_2171__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i22.GSR = "ENABLED";
    FD1S3IX count_2171__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i23.GSR = "ENABLED";
    FD1S3IX count_2171__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i24.GSR = "ENABLED";
    FD1S3IX count_2171__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i25.GSR = "ENABLED";
    FD1S3IX count_2171__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i26.GSR = "ENABLED";
    FD1S3IX count_2171__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i27.GSR = "ENABLED";
    FD1S3IX count_2171__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i28.GSR = "ENABLED";
    FD1S3IX count_2171__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i29.GSR = "ENABLED";
    FD1S3IX count_2171__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i30.GSR = "ENABLED";
    FD1S3IX count_2171__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n28890), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2171__i31.GSR = "ENABLED";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24299), .COUT(n24300), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24298), .COUT(n24299), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24297), .COUT(n24298), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24296), .COUT(n24297), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24295), .COUT(n24296), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24294), .COUT(n24295), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24293), .COUT(n24294), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24293), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1725_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n23961));
    defparam sub_1725_add_2_1.INIT0 = 16'h0000;
    defparam sub_1725_add_2_1.INIT1 = 16'h5999;
    defparam sub_1725_add_2_1.INJECT1_0 = "NO";
    defparam sub_1725_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n28890), .CD(n14388), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_1725_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23970), .COUT(n23971));
    defparam sub_1725_add_2_21.INIT0 = 16'h5999;
    defparam sub_1725_add_2_21.INIT1 = 16'h5999;
    defparam sub_1725_add_2_21.INJECT1_0 = "NO";
    defparam sub_1725_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1725_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23963), .COUT(n23964));
    defparam sub_1725_add_2_7.INIT0 = 16'h5999;
    defparam sub_1725_add_2_7.INIT1 = 16'h5999;
    defparam sub_1725_add_2_7.INJECT1_0 = "NO";
    defparam sub_1725_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1725_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23969), .COUT(n23970));
    defparam sub_1725_add_2_19.INIT0 = 16'h5999;
    defparam sub_1725_add_2_19.INIT1 = 16'h5999;
    defparam sub_1725_add_2_19.INJECT1_0 = "NO";
    defparam sub_1725_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1725_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23968), .COUT(n23969));
    defparam sub_1725_add_2_17.INIT0 = 16'h5999;
    defparam sub_1725_add_2_17.INIT1 = 16'h5999;
    defparam sub_1725_add_2_17.INJECT1_0 = "NO";
    defparam sub_1725_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1725_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23967), .COUT(n23968));
    defparam sub_1725_add_2_15.INIT0 = 16'h5999;
    defparam sub_1725_add_2_15.INIT1 = 16'h5999;
    defparam sub_1725_add_2_15.INJECT1_0 = "NO";
    defparam sub_1725_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24268), .S1(n7156));
    defparam sub_1727_add_2_33.INIT0 = 16'h5999;
    defparam sub_1727_add_2_33.INIT1 = 16'h0000;
    defparam sub_1727_add_2_33.INJECT1_0 = "NO";
    defparam sub_1727_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24267), .COUT(n24268));
    defparam sub_1727_add_2_31.INIT0 = 16'h5999;
    defparam sub_1727_add_2_31.INIT1 = 16'h5999;
    defparam sub_1727_add_2_31.INJECT1_0 = "NO";
    defparam sub_1727_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1725_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n23966), .COUT(n23967));
    defparam sub_1725_add_2_13.INIT0 = 16'h5999;
    defparam sub_1725_add_2_13.INIT1 = 16'h5999;
    defparam sub_1725_add_2_13.INJECT1_0 = "NO";
    defparam sub_1725_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24266), .COUT(n24267));
    defparam sub_1727_add_2_29.INIT0 = 16'h5999;
    defparam sub_1727_add_2_29.INIT1 = 16'h5999;
    defparam sub_1727_add_2_29.INJECT1_0 = "NO";
    defparam sub_1727_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1725_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23976), .S1(n7121));
    defparam sub_1725_add_2_33.INIT0 = 16'h5555;
    defparam sub_1725_add_2_33.INIT1 = 16'h0000;
    defparam sub_1725_add_2_33.INJECT1_0 = "NO";
    defparam sub_1725_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24265), .COUT(n24266));
    defparam sub_1727_add_2_27.INIT0 = 16'h5999;
    defparam sub_1727_add_2_27.INIT1 = 16'h5999;
    defparam sub_1727_add_2_27.INJECT1_0 = "NO";
    defparam sub_1727_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24264), .COUT(n24265));
    defparam sub_1727_add_2_25.INIT0 = 16'h5999;
    defparam sub_1727_add_2_25.INIT1 = 16'h5999;
    defparam sub_1727_add_2_25.INJECT1_0 = "NO";
    defparam sub_1727_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24263), .COUT(n24264));
    defparam sub_1727_add_2_23.INIT0 = 16'h5999;
    defparam sub_1727_add_2_23.INIT1 = 16'h5999;
    defparam sub_1727_add_2_23.INJECT1_0 = "NO";
    defparam sub_1727_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24262), .COUT(n24263));
    defparam sub_1727_add_2_21.INIT0 = 16'h5999;
    defparam sub_1727_add_2_21.INIT1 = 16'h5999;
    defparam sub_1727_add_2_21.INJECT1_0 = "NO";
    defparam sub_1727_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24261), .COUT(n24262));
    defparam sub_1727_add_2_19.INIT0 = 16'h5999;
    defparam sub_1727_add_2_19.INIT1 = 16'h5999;
    defparam sub_1727_add_2_19.INJECT1_0 = "NO";
    defparam sub_1727_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24260), .COUT(n24261));
    defparam sub_1727_add_2_17.INIT0 = 16'h5999;
    defparam sub_1727_add_2_17.INIT1 = 16'h5999;
    defparam sub_1727_add_2_17.INJECT1_0 = "NO";
    defparam sub_1727_add_2_17.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0100000) 
//

module \ArmPeripheral(axis_haddr=8'b0100000)  (read_value, debug_c_c, n11947, 
            GND_net, n30647, n28965, \register_addr[4] , n28899, \register_addr[5] , 
            limit_c_2, n7844, n14, \register_addr[0] , n15, \register_addr[1] , 
            VCC_net, Stepper_Z_nFault_c, n30649, \read_size[0] , n84, 
            Stepper_Z_M0_c_0, n580, prev_select, n28937, n30650, databus, 
            n609, n611, \control_reg[7] , n574, Stepper_Z_Dir_c, Stepper_Z_M2_c_2, 
            Stepper_Z_M1_c_1, \read_size[2] , n60, n30652, n30651, 
            \steps_reg[5] , \steps_reg[3] , n29056, prev_select_adj_143, 
            n28973, n12590, n29011, n29025, \register[2][18] , n29008, 
            n27023, \register[2][19] , n27041, \register[2][20] , n27047, 
            stepping, \register[2][21] , n27048, \register[2][22] , 
            n27040, \register[2][23] , n27039, \register[2][24] , n27035, 
            \register[2][25] , n27050, \register[2][26] , n27024, \register[2][27] , 
            n27049, \register[2][28] , n27044, \register[2][29] , n27032, 
            \register[2][30] , n27037, \register[2][31] , n27043, n29021, 
            \register_addr[2] , n28955, n176, Stepper_Z_En_c, Stepper_Z_Step_c, 
            rw, n28956, n7, \register[2][13] , n27027, n30644, n28918, 
            n26939, n27014, \register[2][14] , n27029, n24970, \register[2][15] , 
            n27038, \register[2][16] , n27031, \register[2][4] , n27030, 
            n28990, n11636, n26917, \register[2][5] , n27034, \register[2][17] , 
            n27033, \register[2][6] , n27036, n22447, n27065, \register[2][7] , 
            n27028, \register[2][8] , n27046, \register[2][9] , n27042, 
            \register[2][10] , n27045, \register[2][11] , n27026, \register[2][12] , 
            n27025, n28991) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    input n11947;
    input GND_net;
    input n30647;
    input n28965;
    input \register_addr[4] ;
    input n28899;
    input \register_addr[5] ;
    input limit_c_2;
    input n7844;
    input n14;
    input \register_addr[0] ;
    input n15;
    input \register_addr[1] ;
    input VCC_net;
    input Stepper_Z_nFault_c;
    input n30649;
    output \read_size[0] ;
    input n84;
    output Stepper_Z_M0_c_0;
    input n580;
    output prev_select;
    input n28937;
    input n30650;
    input [31:0]databus;
    input n609;
    input n611;
    output \control_reg[7] ;
    input n574;
    output Stepper_Z_Dir_c;
    output Stepper_Z_M2_c_2;
    output Stepper_Z_M1_c_1;
    output \read_size[2] ;
    input n60;
    input n30652;
    input n30651;
    output \steps_reg[5] ;
    output \steps_reg[3] ;
    input n29056;
    input prev_select_adj_143;
    input n28973;
    output n12590;
    input n29011;
    input n29025;
    input \register[2][18] ;
    input n29008;
    output n27023;
    input \register[2][19] ;
    output n27041;
    input \register[2][20] ;
    output n27047;
    input stepping;
    input \register[2][21] ;
    output n27048;
    input \register[2][22] ;
    output n27040;
    input \register[2][23] ;
    output n27039;
    input \register[2][24] ;
    output n27035;
    input \register[2][25] ;
    output n27050;
    input \register[2][26] ;
    output n27024;
    input \register[2][27] ;
    output n27049;
    input \register[2][28] ;
    output n27044;
    input \register[2][29] ;
    output n27032;
    input \register[2][30] ;
    output n27037;
    input \register[2][31] ;
    output n27043;
    input n29021;
    input \register_addr[2] ;
    output n28955;
    output n176;
    output Stepper_Z_En_c;
    output Stepper_Z_Step_c;
    input rw;
    input n28956;
    output n7;
    input \register[2][13] ;
    output n27027;
    input n30644;
    input n28918;
    input n26939;
    input n27014;
    input \register[2][14] ;
    output n27029;
    output n24970;
    input \register[2][15] ;
    output n27038;
    input \register[2][16] ;
    output n27031;
    input \register[2][4] ;
    output n27030;
    input n28990;
    input n11636;
    output n26917;
    input \register[2][5] ;
    output n27034;
    input \register[2][17] ;
    output n27033;
    input \register[2][6] ;
    output n27036;
    input n22447;
    output n27065;
    input \register[2][7] ;
    output n27028;
    input \register[2][8] ;
    output n27046;
    input \register[2][9] ;
    output n27042;
    input \register[2][10] ;
    output n27045;
    input \register[2][11] ;
    output n27026;
    input \register[2][12] ;
    output n27025;
    input n28991;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n26969, n26970, n26971, n24388;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]n225;
    
    wire n26972, n26973, n24387, n12086, n12338, n183, n24386, 
        n26966, n26974, n26975, n12324, n24385, n26976, n24384, 
        n18825, n18827, n26977, n24383, n24382, n24381, n26978, 
        n18828;
    wire [31:0]n5778;
    
    wire n26979;
    wire [7:0]n7330;
    
    wire n5, n6, fault_latched;
    wire [31:0]n3273;
    
    wire n24380, prev_step_clk, step_clk, limit_latched, prev_limit_latched;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n24379, n24378, n26980, n26981, n26982, n26983, n26984, 
        n26985, n26986, n26987, n26964, n9600;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n24377, int_step, n20625, n28909, n24376, n24375, n24374, 
        n24373, n26967, n26965, n26968, n27481, n27482, n3272, 
        n49, n62, n58, n50, n27436, n27437, n27438, n41, n60_adj_256, 
        n54, n42, n52, n38, n56, n46;
    wire [31:0]n5742;
    
    wire n27397, n27398, n27399, n27483;
    
    FD1P3AX read_value__i11 (.D(n26969), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n26970), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n26971), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    CCU2D sub_126_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24388), .S0(n225[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_33.INIT0 = 16'h5555;
    defparam sub_126_add_2_33.INIT1 = 16'h0000;
    defparam sub_126_add_2_33.INJECT1_0 = "NO";
    defparam sub_126_add_2_33.INJECT1_1 = "NO";
    FD1P3AX read_value__i14 (.D(n26972), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n26973), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    CCU2D sub_126_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24387), .COUT(n24388), .S0(n225[29]), 
          .S1(n225[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_31.INIT0 = 16'h5555;
    defparam sub_126_add_2_31.INIT1 = 16'h5555;
    defparam sub_126_add_2_31.INJECT1_0 = "NO";
    defparam sub_126_add_2_31.INJECT1_1 = "NO";
    LUT4 i21291_2_lut (.A(n12086), .B(n30647), .Z(n12338)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21291_2_lut.init = 16'heeee;
    LUT4 i21258_4_lut (.A(n28965), .B(\register_addr[4] ), .C(n28899), 
         .D(\register_addr[5] ), .Z(n12086)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i21258_4_lut.init = 16'h1000;
    LUT4 i119_1_lut (.A(limit_c_2), .Z(n183)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i119_1_lut.init = 16'h5555;
    CCU2D sub_126_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24386), .COUT(n24387), .S0(n225[27]), 
          .S1(n225[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_29.INIT0 = 16'h5555;
    defparam sub_126_add_2_29.INIT1 = 16'h5555;
    defparam sub_126_add_2_29.INJECT1_0 = "NO";
    defparam sub_126_add_2_29.INJECT1_1 = "NO";
    FD1P3AX read_value__i16 (.D(n26966), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n26974), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n26975), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(n7844), .B(n30647), .Z(n12324)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    CCU2D sub_126_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24385), .COUT(n24386), .S0(n225[25]), 
          .S1(n225[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_27.INIT0 = 16'h5555;
    defparam sub_126_add_2_27.INIT1 = 16'h5555;
    defparam sub_126_add_2_27.INJECT1_0 = "NO";
    defparam sub_126_add_2_27.INJECT1_1 = "NO";
    FD1P3AX read_value__i19 (.D(n26976), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    CCU2D sub_126_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24384), .COUT(n24385), .S0(n225[23]), 
          .S1(n225[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_25.INIT0 = 16'h5555;
    defparam sub_126_add_2_25.INIT1 = 16'h5555;
    defparam sub_126_add_2_25.INJECT1_0 = "NO";
    defparam sub_126_add_2_25.INJECT1_1 = "NO";
    PFUMX i13085 (.BLUT(n18825), .ALUT(n14), .C0(\register_addr[0] ), 
          .Z(n18827));
    FD1P3AX read_value__i20 (.D(n26977), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    CCU2D sub_126_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24383), .COUT(n24384), .S0(n225[21]), 
          .S1(n225[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_23.INIT0 = 16'h5555;
    defparam sub_126_add_2_23.INIT1 = 16'h5555;
    defparam sub_126_add_2_23.INJECT1_0 = "NO";
    defparam sub_126_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24382), .COUT(n24383), .S0(n225[19]), 
          .S1(n225[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_21.INIT0 = 16'h5555;
    defparam sub_126_add_2_21.INIT1 = 16'h5555;
    defparam sub_126_add_2_21.INJECT1_0 = "NO";
    defparam sub_126_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24381), .COUT(n24382), .S0(n225[17]), 
          .S1(n225[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_19.INIT0 = 16'h5555;
    defparam sub_126_add_2_19.INIT1 = 16'h5555;
    defparam sub_126_add_2_19.INJECT1_0 = "NO";
    defparam sub_126_add_2_19.INJECT1_1 = "NO";
    FD1P3AX read_value__i21 (.D(n26978), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    PFUMX i13088 (.BLUT(n18828), .ALUT(n15), .C0(\register_addr[0] ), 
          .Z(n5778[3]));
    FD1P3AX read_value__i22 (.D(n26979), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    PFUMX i6 (.BLUT(n7330[6]), .ALUT(n5), .C0(\register_addr[1] ), .Z(n6));
    IFS1P3DX fault_latched_179 (.D(Stepper_Z_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_179.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3273[0]), .CK(debug_c_c), .CD(n30649), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n84), .SP(n11947), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    CCU2D sub_126_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24380), .COUT(n24381), .S0(n225[15]), 
          .S1(n225[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_17.INIT0 = 16'h5555;
    defparam sub_126_add_2_17.INIT1 = 16'h5555;
    defparam sub_126_add_2_17.INJECT1_0 = "NO";
    defparam sub_126_add_2_17.INJECT1_1 = "NO";
    FD1P3AX control_reg_i1 (.D(n580), .SP(n12338), .CK(debug_c_c), .Q(Stepper_Z_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_176 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_176.GSR = "ENABLED";
    FD1S3AX limit_latched_177 (.D(n183), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_177.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_178 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_178.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n580), .SP(n12324), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_175 (.D(n28937), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_175.GSR = "ENABLED";
    CCU2D sub_126_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24379), .COUT(n24380), .S0(n225[13]), 
          .S1(n225[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_15.INIT0 = 16'h5555;
    defparam sub_126_add_2_15.INIT1 = 16'h5555;
    defparam sub_126_add_2_15.INJECT1_0 = "NO";
    defparam sub_126_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24378), .COUT(n24379), .S0(n225[11]), 
          .S1(n225[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_13.INIT0 = 16'h5555;
    defparam sub_126_add_2_13.INIT1 = 16'h5555;
    defparam sub_126_add_2_13.INJECT1_0 = "NO";
    defparam sub_126_add_2_13.INJECT1_1 = "NO";
    FD1P3AX read_value__i23 (.D(n26980), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n26981), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n26982), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n26983), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n26984), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n26985), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n26986), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n26987), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n26964), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n7844), .PD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n7844), .PD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n7844), .PD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n7844), .PD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n7844), .PD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n7844), .PD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n7844), .PD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n609), .SP(n12324), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n611), .SP(n12324), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n12086), .CD(n9600), .CK(debug_c_c), 
            .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3AX control_reg_i7 (.D(n574), .SP(n12338), .CK(debug_c_c), .Q(control_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n12086), .PD(n30650), 
            .CK(debug_c_c), .Q(Stepper_Z_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n609), .SP(n12338), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n12086), .PD(n30650), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n611), .SP(n12338), .CK(debug_c_c), .Q(Stepper_Z_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n12086), .PD(n30650), 
            .CK(debug_c_c), .Q(Stepper_Z_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    CCU2D sub_126_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24377), .COUT(n24378), .S0(n225[9]), .S1(n225[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_11.INIT0 = 16'h5555;
    defparam sub_126_add_2_11.INIT1 = 16'h5555;
    defparam sub_126_add_2_11.INJECT1_0 = "NO";
    defparam sub_126_add_2_11.INJECT1_1 = "NO";
    FD1P3AX int_step_183 (.D(n28909), .SP(n20625), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_183.GSR = "ENABLED";
    CCU2D sub_126_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24376), .COUT(n24377), .S0(n225[7]), .S1(n225[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_9.INIT0 = 16'h5555;
    defparam sub_126_add_2_9.INIT1 = 16'h5555;
    defparam sub_126_add_2_9.INJECT1_0 = "NO";
    defparam sub_126_add_2_9.INJECT1_1 = "NO";
    FD1P3AX read_size__i2 (.D(n60), .SP(n11947), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3273[31]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3273[30]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3273[29]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3273[28]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3273[27]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3273[26]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3273[25]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3273[24]), .CK(debug_c_c), .CD(n30652), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3273[23]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3273[22]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3273[21]), .CK(debug_c_c), .CD(n30650), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3273[20]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3273[19]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3273[18]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3273[17]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3273[16]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3273[15]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3273[14]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3273[13]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3273[12]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3273[11]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3273[10]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3273[9]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3273[8]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3273[7]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3273[6]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3273[5]), .CK(debug_c_c), .CD(n30651), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3273[4]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3273[3]), .CK(debug_c_c), .CD(n30651), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3273[2]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3273[1]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    CCU2D sub_126_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24375), .COUT(n24376), .S0(n225[5]), .S1(n225[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_7.INIT0 = 16'h5555;
    defparam sub_126_add_2_7.INIT1 = 16'h5555;
    defparam sub_126_add_2_7.INJECT1_0 = "NO";
    defparam sub_126_add_2_7.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(n29056), .B(n30647), .C(prev_select_adj_143), .D(n28973), 
         .Z(n12590)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n29011), .B(n29025), .C(\register[2][18] ), 
         .D(n29008), .Z(n27023)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    CCU2D sub_126_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24374), .COUT(n24375), .S0(n225[3]), .S1(n225[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_5.INIT0 = 16'h5555;
    defparam sub_126_add_2_5.INIT1 = 16'h5555;
    defparam sub_126_add_2_5.INJECT1_0 = "NO";
    defparam sub_126_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24373), .COUT(n24374), .S0(n225[1]), .S1(n225[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_3.INIT0 = 16'h5555;
    defparam sub_126_add_2_3.INIT1 = 16'h5555;
    defparam sub_126_add_2_3.INJECT1_0 = "NO";
    defparam sub_126_add_2_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_188 (.A(n29011), .B(n29025), .C(\register[2][19] ), 
         .D(n29008), .Z(n27041)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_188.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_189 (.A(n29011), .B(n29025), .C(\register[2][20] ), 
         .D(n29008), .Z(n27047)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_189.init = 16'h1000;
    CCU2D sub_126_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(stepping), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n24373), .S1(n225[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_1.INIT0 = 16'h0000;
    defparam sub_126_add_2_1.INIT1 = 16'h5595;
    defparam sub_126_add_2_1.INJECT1_0 = "NO";
    defparam sub_126_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_190 (.A(n29011), .B(n29025), .C(\register[2][21] ), 
         .D(n29008), .Z(n27048)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_190.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_191 (.A(n29011), .B(n29025), .C(\register[2][22] ), 
         .D(n29008), .Z(n27040)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_191.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_192 (.A(n29011), .B(n29025), .C(\register[2][23] ), 
         .D(n29008), .Z(n27039)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_192.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_193 (.A(n29011), .B(n29025), .C(\register[2][24] ), 
         .D(n29008), .Z(n27035)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_193.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_194 (.A(n29011), .B(n29025), .C(\register[2][25] ), 
         .D(n29008), .Z(n27050)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_194.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_195 (.A(n29011), .B(n29025), .C(\register[2][26] ), 
         .D(n29008), .Z(n27024)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_195.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_196 (.A(n29011), .B(n29025), .C(\register[2][27] ), 
         .D(n29008), .Z(n27049)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_196.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_197 (.A(n29011), .B(n29025), .C(\register[2][28] ), 
         .D(n29008), .Z(n27044)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_197.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_198 (.A(n29011), .B(n29025), .C(\register[2][29] ), 
         .D(n29008), .Z(n27032)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_198.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_199 (.A(n29011), .B(n29025), .C(\register[2][30] ), 
         .D(n29008), .Z(n27037)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_199.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_200 (.A(n29011), .B(n29025), .C(\register[2][31] ), 
         .D(n29008), .Z(n27043)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_200.init = 16'h1000;
    LUT4 i1_3_lut_rep_297_4_lut (.A(n29011), .B(n29025), .C(n29021), .D(\register_addr[2] ), 
         .Z(n28955)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_3_lut_rep_297_4_lut.init = 16'hfeee;
    LUT4 i14652_1_lut_3_lut_4_lut (.A(n29011), .B(n29025), .C(n29021), 
         .D(\register_addr[2] ), .Z(n176)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;
    defparam i14652_1_lut_3_lut_4_lut.init = 16'h0111;
    LUT4 i1_4_lut (.A(div_factor_reg[8]), .B(\register_addr[1] ), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n26967)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_201 (.A(div_factor_reg[9]), .B(\register_addr[1] ), 
         .C(steps_reg[9]), .D(\register_addr[0] ), .Z(n26965)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_201.init = 16'hc088;
    LUT4 i2_3_lut_rep_251 (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .Z(n28909)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i2_3_lut_rep_251.init = 16'h0808;
    LUT4 i1_4_lut_adj_202 (.A(div_factor_reg[10]), .B(\register_addr[1] ), 
         .C(steps_reg[10]), .D(\register_addr[0] ), .Z(n26968)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_202.init = 16'hc088;
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    LUT4 i13083_3_lut (.A(Stepper_Z_Dir_c), .B(div_factor_reg[5]), .C(\register_addr[1] ), 
         .Z(n18825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13083_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    LUT4 i14880_4_lut_4_lut (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .D(n30647), .Z(n20625)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i14880_4_lut_4_lut.init = 16'h0038;
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n12324), .CD(n30650), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 i21111_3_lut (.A(Stepper_Z_M2_c_2), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n27481)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21111_3_lut.init = 16'hcaca;
    LUT4 i21112_3_lut (.A(div_factor_reg[2]), .B(steps_reg[2]), .C(\register_addr[0] ), 
         .Z(n27482)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21112_3_lut.init = 16'hcaca;
    LUT4 i8_1_lut (.A(control_reg[6]), .Z(Stepper_Z_En_c)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(44[14:29])
    defparam i8_1_lut.init = 16'h5555;
    LUT4 i21204_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_Z_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i21204_2_lut.init = 16'h9999;
    LUT4 i1_4_lut_adj_203 (.A(div_factor_reg[20]), .B(\register_addr[1] ), 
         .C(steps_reg[20]), .D(\register_addr[0] ), .Z(n26977)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_203.init = 16'hc088;
    LUT4 i1_4_lut_adj_204 (.A(div_factor_reg[11]), .B(\register_addr[1] ), 
         .C(steps_reg[11]), .D(\register_addr[0] ), .Z(n26969)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_204.init = 16'hc088;
    LUT4 i1_4_lut_adj_205 (.A(div_factor_reg[23]), .B(\register_addr[1] ), 
         .C(steps_reg[23]), .D(\register_addr[0] ), .Z(n26980)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_205.init = 16'hc088;
    LUT4 i2_2_lut_4_lut (.A(n28965), .B(\register_addr[4] ), .C(rw), .D(n28956), 
         .Z(n7)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i2_2_lut_4_lut.init = 16'hfffb;
    LUT4 i1_4_lut_adj_206 (.A(div_factor_reg[12]), .B(\register_addr[1] ), 
         .C(steps_reg[12]), .D(\register_addr[0] ), .Z(n26970)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_206.init = 16'hc088;
    LUT4 i1_4_lut_adj_207 (.A(div_factor_reg[13]), .B(\register_addr[1] ), 
         .C(steps_reg[13]), .D(\register_addr[0] ), .Z(n26971)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_207.init = 16'hc088;
    LUT4 i1_4_lut_adj_208 (.A(div_factor_reg[14]), .B(\register_addr[1] ), 
         .C(steps_reg[14]), .D(\register_addr[0] ), .Z(n26972)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_208.init = 16'hc088;
    LUT4 i1_4_lut_adj_209 (.A(div_factor_reg[21]), .B(\register_addr[1] ), 
         .C(steps_reg[21]), .D(\register_addr[0] ), .Z(n26978)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_209.init = 16'hc088;
    LUT4 i13086_3_lut (.A(control_reg[3]), .B(div_factor_reg[3]), .C(\register_addr[1] ), 
         .Z(n18828)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13086_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_210 (.A(div_factor_reg[24]), .B(\register_addr[1] ), 
         .C(steps_reg[24]), .D(\register_addr[0] ), .Z(n26981)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_210.init = 16'hc088;
    LUT4 i1_4_lut_adj_211 (.A(div_factor_reg[25]), .B(\register_addr[1] ), 
         .C(steps_reg[25]), .D(\register_addr[0] ), .Z(n26982)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_211.init = 16'hc088;
    LUT4 i1_4_lut_adj_212 (.A(div_factor_reg[31]), .B(\register_addr[1] ), 
         .C(steps_reg[31]), .D(\register_addr[0] ), .Z(n26964)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_212.init = 16'hc088;
    LUT4 i1_4_lut_adj_213 (.A(div_factor_reg[26]), .B(\register_addr[1] ), 
         .C(steps_reg[26]), .D(\register_addr[0] ), .Z(n26983)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_213.init = 16'hc088;
    LUT4 i1_4_lut_adj_214 (.A(div_factor_reg[27]), .B(\register_addr[1] ), 
         .C(steps_reg[27]), .D(\register_addr[0] ), .Z(n26984)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_214.init = 16'hc088;
    LUT4 i1_4_lut_adj_215 (.A(div_factor_reg[28]), .B(\register_addr[1] ), 
         .C(steps_reg[28]), .D(\register_addr[0] ), .Z(n26985)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_215.init = 16'hc088;
    LUT4 i1_4_lut_adj_216 (.A(div_factor_reg[29]), .B(\register_addr[1] ), 
         .C(steps_reg[29]), .D(\register_addr[0] ), .Z(n26986)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_216.init = 16'hc088;
    LUT4 i1_4_lut_adj_217 (.A(div_factor_reg[30]), .B(\register_addr[1] ), 
         .C(steps_reg[30]), .D(\register_addr[0] ), .Z(n26987)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_217.init = 16'hc088;
    LUT4 i1_2_lut_3_lut_4_lut_adj_218 (.A(n29011), .B(n29025), .C(\register[2][13] ), 
         .D(n29008), .Z(n27027)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_218.init = 16'h1000;
    LUT4 i2_3_lut_4_lut (.A(n30644), .B(n28918), .C(n26939), .D(n27014), 
         .Z(n3272)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i2_3_lut_4_lut.init = 16'h4000;
    LUT4 i3839_3_lut (.A(prev_limit_latched), .B(n30647), .C(limit_latched), 
         .Z(n9600)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i3839_3_lut.init = 16'hdcdc;
    LUT4 i1_2_lut_3_lut_4_lut_adj_219 (.A(n29011), .B(n29025), .C(\register[2][14] ), 
         .D(n29008), .Z(n27029)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_219.init = 16'h1000;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n24970)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    PFUMX i21068 (.BLUT(n27436), .ALUT(n27437), .C0(\register_addr[1] ), 
          .Z(n27438));
    LUT4 i17_4_lut (.A(steps_reg[0]), .B(steps_reg[9]), .C(steps_reg[28]), 
         .D(steps_reg[2]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_220 (.A(div_factor_reg[22]), .B(\register_addr[1] ), 
         .C(steps_reg[22]), .D(\register_addr[0] ), .Z(n26979)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_220.init = 16'hc088;
    LUT4 i30_4_lut (.A(n41), .B(n60_adj_256), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i14105_2_lut (.A(control_reg[6]), .B(\register_addr[0] ), .Z(n7330[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14105_2_lut.init = 16'h2222;
    LUT4 i5_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i5_3_lut.init = 16'hcaca;
    LUT4 i21066_3_lut (.A(Stepper_Z_M0_c_0), .B(stepping), .C(\register_addr[0] ), 
         .Z(n27436)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21066_3_lut.init = 16'hcaca;
    LUT4 i21067_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n27437)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21067_3_lut.init = 16'hcaca;
    LUT4 i26_4_lut (.A(steps_reg[25]), .B(n52), .C(n38), .D(steps_reg[26]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_221 (.A(div_factor_reg[19]), .B(\register_addr[1] ), 
         .C(steps_reg[19]), .D(\register_addr[0] ), .Z(n26976)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_221.init = 16'hc088;
    LUT4 i14106_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n7330[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14106_2_lut.init = 16'h2222;
    LUT4 i18_4_lut (.A(steps_reg[8]), .B(steps_reg[11]), .C(steps_reg[16]), 
         .D(steps_reg[21]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[30]), .B(steps_reg[7]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[20]), .B(n56), .C(n46), .D(steps_reg[15]), 
         .Z(n60_adj_256)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[22]), .B(steps_reg[12]), .C(steps_reg[6]), 
         .D(steps_reg[18]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[14]), .B(steps_reg[19]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[13]), .B(steps_reg[17]), .C(\steps_reg[5] ), 
         .D(steps_reg[31]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[23]), .B(steps_reg[29]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[27]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[10]), .B(\steps_reg[3] ), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 mux_1642_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n5742[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1642_i5_3_lut.init = 16'hcaca;
    LUT4 i14104_2_lut (.A(\control_reg[7] ), .B(\register_addr[0] ), .Z(n7330[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14104_2_lut.init = 16'h2222;
    LUT4 mux_1334_i1_3_lut (.A(n225[0]), .B(databus[0]), .C(n3272), .Z(n3273[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n5742[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1642_i8_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_222 (.A(n29011), .B(n29025), .C(\register[2][15] ), 
         .D(n29008), .Z(n27038)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_222.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_223 (.A(n29011), .B(n29025), .C(\register[2][16] ), 
         .D(n29008), .Z(n27031)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_223.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_224 (.A(n29011), .B(n29025), .C(\register[2][4] ), 
         .D(n29008), .Z(n27030)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_224.init = 16'h1000;
    LUT4 i1_4_lut_adj_225 (.A(div_factor_reg[15]), .B(\register_addr[1] ), 
         .C(steps_reg[15]), .D(\register_addr[0] ), .Z(n26973)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_225.init = 16'hc088;
    LUT4 i1_4_lut_adj_226 (.A(div_factor_reg[16]), .B(\register_addr[1] ), 
         .C(steps_reg[16]), .D(\register_addr[0] ), .Z(n26966)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_226.init = 16'hc088;
    LUT4 i1_4_lut_adj_227 (.A(div_factor_reg[17]), .B(\register_addr[1] ), 
         .C(steps_reg[17]), .D(\register_addr[0] ), .Z(n26974)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_227.init = 16'hc088;
    LUT4 i1_4_lut_adj_228 (.A(div_factor_reg[18]), .B(\register_addr[1] ), 
         .C(steps_reg[18]), .D(\register_addr[0] ), .Z(n26975)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_228.init = 16'hc088;
    LUT4 i1_2_lut_3_lut_4_lut_adj_229 (.A(n28990), .B(n11636), .C(\register_addr[1] ), 
         .D(n12590), .Z(n26917)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C)+!B !((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_3_lut_4_lut_adj_229.init = 16'h40f0;
    LUT4 mux_1334_i32_3_lut (.A(n225[31]), .B(databus[31]), .C(n3272), 
         .Z(n3273[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i31_3_lut (.A(n225[30]), .B(databus[30]), .C(n3272), 
         .Z(n3273[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i30_3_lut (.A(n225[29]), .B(databus[29]), .C(n3272), 
         .Z(n3273[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i29_3_lut (.A(n225[28]), .B(databus[28]), .C(n3272), 
         .Z(n3273[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i28_3_lut (.A(n225[27]), .B(databus[27]), .C(n3272), 
         .Z(n3273[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i27_3_lut (.A(n225[26]), .B(databus[26]), .C(n3272), 
         .Z(n3273[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i26_3_lut (.A(n225[25]), .B(databus[25]), .C(n3272), 
         .Z(n3273[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i25_3_lut (.A(n225[24]), .B(databus[24]), .C(n3272), 
         .Z(n3273[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i24_3_lut (.A(n225[23]), .B(databus[23]), .C(n3272), 
         .Z(n3273[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i23_3_lut (.A(n225[22]), .B(databus[22]), .C(n3272), 
         .Z(n3273[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i22_3_lut (.A(n225[21]), .B(databus[21]), .C(n3272), 
         .Z(n3273[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i21_3_lut (.A(n225[20]), .B(databus[20]), .C(n3272), 
         .Z(n3273[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i20_3_lut (.A(n225[19]), .B(databus[19]), .C(n3272), 
         .Z(n3273[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i19_3_lut (.A(n225[18]), .B(databus[18]), .C(n3272), 
         .Z(n3273[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i18_3_lut (.A(n225[17]), .B(databus[17]), .C(n3272), 
         .Z(n3273[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i17_3_lut (.A(n225[16]), .B(databus[16]), .C(n3272), 
         .Z(n3273[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i16_3_lut (.A(n225[15]), .B(databus[15]), .C(n3272), 
         .Z(n3273[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i16_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i0 (.D(n27438), .SP(n11947), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 mux_1334_i15_3_lut (.A(n225[14]), .B(databus[14]), .C(n3272), 
         .Z(n3273[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i15_3_lut.init = 16'hcaca;
    PFUMX i21029 (.BLUT(n27397), .ALUT(n27398), .C0(\register_addr[1] ), 
          .Z(n27399));
    LUT4 mux_1334_i14_3_lut (.A(n225[13]), .B(databus[13]), .C(n3272), 
         .Z(n3273[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i13_3_lut (.A(n225[12]), .B(databus[12]), .C(n3272), 
         .Z(n3273[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i12_3_lut (.A(n225[11]), .B(databus[11]), .C(n3272), 
         .Z(n3273[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i12_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_230 (.A(n29011), .B(n29025), .C(\register[2][5] ), 
         .D(n29008), .Z(n27034)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_230.init = 16'h1000;
    PFUMX mux_1646_i5 (.BLUT(n7330[4]), .ALUT(n5742[4]), .C0(\register_addr[1] ), 
          .Z(n5778[4]));
    PFUMX mux_1646_i8 (.BLUT(n7330[7]), .ALUT(n5742[7]), .C0(\register_addr[1] ), 
          .Z(n5778[7]));
    LUT4 mux_1334_i11_3_lut (.A(n225[10]), .B(databus[10]), .C(n3272), 
         .Z(n3273[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i10_3_lut (.A(n225[9]), .B(databus[9]), .C(n3272), .Z(n3273[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i9_3_lut (.A(n225[8]), .B(databus[8]), .C(n3272), .Z(n3273[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i9_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_231 (.A(n29011), .B(n29025), .C(\register[2][17] ), 
         .D(n29008), .Z(n27033)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_231.init = 16'h1000;
    LUT4 mux_1334_i8_3_lut (.A(n225[7]), .B(databus[7]), .C(n3272), .Z(n3273[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i8_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i1 (.D(n27399), .SP(n11947), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n27483), .SP(n11947), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n5778[3]), .SP(n11947), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    LUT4 mux_1334_i7_3_lut (.A(n225[6]), .B(databus[6]), .C(n3272), .Z(n3273[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i7_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i4 (.D(n5778[4]), .SP(n11947), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    LUT4 mux_1334_i6_3_lut (.A(n225[5]), .B(databus[5]), .C(n3272), .Z(n3273[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1334_i5_3_lut (.A(n225[4]), .B(databus[4]), .C(n3272), .Z(n3273[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i5_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i5 (.D(n18827), .SP(n11947), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6), .SP(n11947), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    LUT4 mux_1334_i4_3_lut (.A(n225[3]), .B(databus[3]), .C(n3272), .Z(n3273[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i4_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i7 (.D(n5778[7]), .SP(n11947), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_232 (.A(n29011), .B(n29025), .C(\register[2][6] ), 
         .D(n29008), .Z(n27036)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_232.init = 16'h1000;
    LUT4 mux_1334_i3_3_lut (.A(n225[2]), .B(databus[2]), .C(n3272), .Z(n3273[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i3_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i8 (.D(n26967), .SP(n11947), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n26965), .SP(n11947), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    LUT4 mux_1334_i2_3_lut (.A(n225[1]), .B(databus[1]), .C(n3272), .Z(n3273[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1334_i2_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i10 (.D(n26968), .SP(n11947), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    LUT4 i21277_3_lut_4_lut (.A(n29011), .B(n29025), .C(\register_addr[2] ), 
         .D(n22447), .Z(n27065)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;
    defparam i21277_3_lut_4_lut.init = 16'h0111;
    LUT4 i1_2_lut_3_lut_4_lut_adj_233 (.A(n29011), .B(n29025), .C(\register[2][7] ), 
         .D(n29008), .Z(n27028)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_233.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_234 (.A(n29011), .B(n29025), .C(\register[2][8] ), 
         .D(n29008), .Z(n27046)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_234.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_235 (.A(n29011), .B(n29025), .C(\register[2][9] ), 
         .D(n29008), .Z(n27042)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_235.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_236 (.A(n29011), .B(n29025), .C(\register[2][10] ), 
         .D(n29008), .Z(n27045)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_236.init = 16'h1000;
    LUT4 i21027_3_lut (.A(Stepper_Z_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n27397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21027_3_lut.init = 16'hcaca;
    LUT4 i21028_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n27398)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21028_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_237 (.A(n29011), .B(n29025), .C(\register[2][11] ), 
         .D(n29008), .Z(n27026)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_237.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_238 (.A(n29011), .B(n29025), .C(\register[2][12] ), 
         .D(n29008), .Z(n27025)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_238.init = 16'h1000;
    PFUMX i21113 (.BLUT(n27481), .ALUT(n27482), .C0(\register_addr[1] ), 
          .Z(n27483));
    ClockDivider step_clk_gen (.GND_net(GND_net), .step_clk(step_clk), .debug_c_c(debug_c_c), 
            .n28991(n28991), .n30647(n30647), .div_factor_reg({div_factor_reg})) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider
//

module ClockDivider (GND_net, step_clk, debug_c_c, n28991, n30647, 
            div_factor_reg) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output step_clk;
    input debug_c_c;
    input n28991;
    input n30647;
    input [31:0]div_factor_reg;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n24063;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n24064, n24062, n24061, n24060, n24059, n24058, n24057, 
        n7017, n24056;
    wire [31:0]n40;
    
    wire n7052, n24055, n28891;
    wire [31:0]n134;
    
    wire n24054, n24053, n7086, n14373, n24052, n24051, n24050, 
        n24049, n24459, n24458, n24457, n24324, n24323, n24456, 
        n24455, n24048, n24322, n24321, n24454, n24047, n24320, 
        n24453, n24046, n24452, n24451, n24450, n24319, n24318, 
        n24449, n24448, n24317, n24447, n24316, n24446, n24315, 
        n24045, n24445, n24444, n24314, n24313, n24312, n24311, 
        n24310, n24309, n24044, n24043, n24042, n24041, n24040, 
        n24039, n24038, n24037, n24036, n24035, n24034, n24033, 
        n24032, n24031, n24030, n24029, n24028, n24027, n24026, 
        n24025, n24072, n24071, n24070, n24069, n24068, n24067, 
        n24066, n24065;
    
    CCU2D sub_1720_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24063), .COUT(n24064));
    defparam sub_1720_add_2_15.INIT0 = 16'h5999;
    defparam sub_1720_add_2_15.INIT1 = 16'h5999;
    defparam sub_1720_add_2_15.INJECT1_0 = "NO";
    defparam sub_1720_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1720_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24062), .COUT(n24063));
    defparam sub_1720_add_2_13.INIT0 = 16'h5999;
    defparam sub_1720_add_2_13.INIT1 = 16'h5999;
    defparam sub_1720_add_2_13.INJECT1_0 = "NO";
    defparam sub_1720_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1720_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24061), .COUT(n24062));
    defparam sub_1720_add_2_11.INIT0 = 16'h5999;
    defparam sub_1720_add_2_11.INIT1 = 16'h5999;
    defparam sub_1720_add_2_11.INJECT1_0 = "NO";
    defparam sub_1720_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1720_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24060), .COUT(n24061));
    defparam sub_1720_add_2_9.INIT0 = 16'h5999;
    defparam sub_1720_add_2_9.INIT1 = 16'h5999;
    defparam sub_1720_add_2_9.INJECT1_0 = "NO";
    defparam sub_1720_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1720_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24059), .COUT(n24060));
    defparam sub_1720_add_2_7.INIT0 = 16'h5999;
    defparam sub_1720_add_2_7.INIT1 = 16'h5999;
    defparam sub_1720_add_2_7.INJECT1_0 = "NO";
    defparam sub_1720_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1720_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24058), .COUT(n24059));
    defparam sub_1720_add_2_5.INIT0 = 16'h5999;
    defparam sub_1720_add_2_5.INIT1 = 16'h5999;
    defparam sub_1720_add_2_5.INJECT1_0 = "NO";
    defparam sub_1720_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1720_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24057), .COUT(n24058));
    defparam sub_1720_add_2_3.INIT0 = 16'h5999;
    defparam sub_1720_add_2_3.INIT1 = 16'h5999;
    defparam sub_1720_add_2_3.INJECT1_0 = "NO";
    defparam sub_1720_add_2_3.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n7017), .CK(debug_c_c), .CD(n28991), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_1720_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n24057));
    defparam sub_1720_add_2_1.INIT0 = 16'h0000;
    defparam sub_1720_add_2_1.INIT1 = 16'h5999;
    defparam sub_1720_add_2_1.INJECT1_0 = "NO";
    defparam sub_1720_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24056), .S1(n7052));
    defparam sub_1722_add_2_33.INIT0 = 16'h5999;
    defparam sub_1722_add_2_33.INIT1 = 16'h0000;
    defparam sub_1722_add_2_33.INJECT1_0 = "NO";
    defparam sub_1722_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24055), .COUT(n24056));
    defparam sub_1722_add_2_31.INIT0 = 16'h5999;
    defparam sub_1722_add_2_31.INIT1 = 16'h5999;
    defparam sub_1722_add_2_31.INJECT1_0 = "NO";
    defparam sub_1722_add_2_31.INJECT1_1 = "NO";
    FD1S3IX count_2170__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i0.GSR = "ENABLED";
    LUT4 i958_2_lut_rep_233 (.A(n7052), .B(n30647), .Z(n28891)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i958_2_lut_rep_233.init = 16'heeee;
    CCU2D sub_1722_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24054), .COUT(n24055));
    defparam sub_1722_add_2_29.INIT0 = 16'h5999;
    defparam sub_1722_add_2_29.INIT1 = 16'h5999;
    defparam sub_1722_add_2_29.INJECT1_0 = "NO";
    defparam sub_1722_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24053), .COUT(n24054));
    defparam sub_1722_add_2_27.INIT0 = 16'h5999;
    defparam sub_1722_add_2_27.INIT1 = 16'h5999;
    defparam sub_1722_add_2_27.INJECT1_0 = "NO";
    defparam sub_1722_add_2_27.INJECT1_1 = "NO";
    LUT4 i8607_2_lut_3_lut (.A(n7052), .B(n30647), .C(n7086), .Z(n14373)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i8607_2_lut_3_lut.init = 16'he0e0;
    CCU2D sub_1722_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24052), .COUT(n24053));
    defparam sub_1722_add_2_25.INIT0 = 16'h5999;
    defparam sub_1722_add_2_25.INIT1 = 16'h5999;
    defparam sub_1722_add_2_25.INJECT1_0 = "NO";
    defparam sub_1722_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24051), .COUT(n24052));
    defparam sub_1722_add_2_23.INIT0 = 16'h5999;
    defparam sub_1722_add_2_23.INIT1 = 16'h5999;
    defparam sub_1722_add_2_23.INJECT1_0 = "NO";
    defparam sub_1722_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24050), .COUT(n24051));
    defparam sub_1722_add_2_21.INIT0 = 16'h5999;
    defparam sub_1722_add_2_21.INIT1 = 16'h5999;
    defparam sub_1722_add_2_21.INJECT1_0 = "NO";
    defparam sub_1722_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24049), .COUT(n24050));
    defparam sub_1722_add_2_19.INIT0 = 16'h5999;
    defparam sub_1722_add_2_19.INIT1 = 16'h5999;
    defparam sub_1722_add_2_19.INJECT1_0 = "NO";
    defparam sub_1722_add_2_19.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    CCU2D count_2170_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24459), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_33.INIT1 = 16'h0000;
    defparam count_2170_add_4_33.INJECT1_0 = "NO";
    defparam count_2170_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24458), .COUT(n24459), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2170_add_4_31.INJECT1_0 = "NO";
    defparam count_2170_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24457), .COUT(n24458), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2170_add_4_29.INJECT1_0 = "NO";
    defparam count_2170_add_4_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24324), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24323), .COUT(n24324), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24456), .COUT(n24457), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2170_add_4_27.INJECT1_0 = "NO";
    defparam count_2170_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24455), .COUT(n24456), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2170_add_4_25.INJECT1_0 = "NO";
    defparam count_2170_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24048), .COUT(n24049));
    defparam sub_1722_add_2_17.INIT0 = 16'h5999;
    defparam sub_1722_add_2_17.INIT1 = 16'h5999;
    defparam sub_1722_add_2_17.INJECT1_0 = "NO";
    defparam sub_1722_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24322), .COUT(n24323), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24321), .COUT(n24322), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24454), .COUT(n24455), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2170_add_4_23.INJECT1_0 = "NO";
    defparam count_2170_add_4_23.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24047), .COUT(n24048));
    defparam sub_1722_add_2_15.INIT0 = 16'h5999;
    defparam sub_1722_add_2_15.INIT1 = 16'h5999;
    defparam sub_1722_add_2_15.INJECT1_0 = "NO";
    defparam sub_1722_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24320), .COUT(n24321), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24453), .COUT(n24454), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2170_add_4_21.INJECT1_0 = "NO";
    defparam count_2170_add_4_21.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24046), .COUT(n24047));
    defparam sub_1722_add_2_13.INIT0 = 16'h5999;
    defparam sub_1722_add_2_13.INIT1 = 16'h5999;
    defparam sub_1722_add_2_13.INJECT1_0 = "NO";
    defparam sub_1722_add_2_13.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24452), .COUT(n24453), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2170_add_4_19.INJECT1_0 = "NO";
    defparam count_2170_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24451), .COUT(n24452), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2170_add_4_17.INJECT1_0 = "NO";
    defparam count_2170_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24450), .COUT(n24451), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2170_add_4_15.INJECT1_0 = "NO";
    defparam count_2170_add_4_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24319), .COUT(n24320), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24318), .COUT(n24319), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24449), .COUT(n24450), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2170_add_4_13.INJECT1_0 = "NO";
    defparam count_2170_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24448), .COUT(n24449), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2170_add_4_11.INJECT1_0 = "NO";
    defparam count_2170_add_4_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24317), .COUT(n24318), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24447), .COUT(n24448), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2170_add_4_9.INJECT1_0 = "NO";
    defparam count_2170_add_4_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24316), .COUT(n24317), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24446), .COUT(n24447), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2170_add_4_7.INJECT1_0 = "NO";
    defparam count_2170_add_4_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24315), .COUT(n24316), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24045), .COUT(n24046));
    defparam sub_1722_add_2_11.INIT0 = 16'h5999;
    defparam sub_1722_add_2_11.INIT1 = 16'h5999;
    defparam sub_1722_add_2_11.INJECT1_0 = "NO";
    defparam sub_1722_add_2_11.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24445), .COUT(n24446), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2170_add_4_5.INJECT1_0 = "NO";
    defparam count_2170_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24444), .COUT(n24445), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2170_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2170_add_4_3.INJECT1_0 = "NO";
    defparam count_2170_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2170_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24444), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170_add_4_1.INIT0 = 16'hF000;
    defparam count_2170_add_4_1.INIT1 = 16'h0555;
    defparam count_2170_add_4_1.INJECT1_0 = "NO";
    defparam count_2170_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24314), .COUT(n24315), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24313), .COUT(n24314), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n28891), .PD(n14373), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24312), .COUT(n24313), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24311), .COUT(n24312), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24310), .COUT(n24311), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24309), .COUT(n24310), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24309), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24044), .COUT(n24045));
    defparam sub_1722_add_2_9.INIT0 = 16'h5999;
    defparam sub_1722_add_2_9.INIT1 = 16'h5999;
    defparam sub_1722_add_2_9.INJECT1_0 = "NO";
    defparam sub_1722_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24043), .COUT(n24044));
    defparam sub_1722_add_2_7.INIT0 = 16'h5999;
    defparam sub_1722_add_2_7.INIT1 = 16'h5999;
    defparam sub_1722_add_2_7.INJECT1_0 = "NO";
    defparam sub_1722_add_2_7.INJECT1_1 = "NO";
    FD1S3IX count_2170__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i1.GSR = "ENABLED";
    CCU2D sub_1722_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24042), .COUT(n24043));
    defparam sub_1722_add_2_5.INIT0 = 16'h5999;
    defparam sub_1722_add_2_5.INIT1 = 16'h5999;
    defparam sub_1722_add_2_5.INJECT1_0 = "NO";
    defparam sub_1722_add_2_5.INJECT1_1 = "NO";
    FD1S3IX count_2170__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i2.GSR = "ENABLED";
    FD1S3IX count_2170__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i3.GSR = "ENABLED";
    FD1S3IX count_2170__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i4.GSR = "ENABLED";
    FD1S3IX count_2170__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i5.GSR = "ENABLED";
    FD1S3IX count_2170__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i6.GSR = "ENABLED";
    FD1S3IX count_2170__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i7.GSR = "ENABLED";
    FD1S3IX count_2170__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i8.GSR = "ENABLED";
    FD1S3IX count_2170__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i9.GSR = "ENABLED";
    FD1S3IX count_2170__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i10.GSR = "ENABLED";
    FD1S3IX count_2170__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i11.GSR = "ENABLED";
    FD1S3IX count_2170__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i12.GSR = "ENABLED";
    FD1S3IX count_2170__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i13.GSR = "ENABLED";
    FD1S3IX count_2170__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i14.GSR = "ENABLED";
    FD1S3IX count_2170__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i15.GSR = "ENABLED";
    FD1S3IX count_2170__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i16.GSR = "ENABLED";
    FD1S3IX count_2170__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i17.GSR = "ENABLED";
    FD1S3IX count_2170__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i18.GSR = "ENABLED";
    FD1S3IX count_2170__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i19.GSR = "ENABLED";
    FD1S3IX count_2170__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i20.GSR = "ENABLED";
    FD1S3IX count_2170__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i21.GSR = "ENABLED";
    FD1S3IX count_2170__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i22.GSR = "ENABLED";
    FD1S3IX count_2170__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i23.GSR = "ENABLED";
    FD1S3IX count_2170__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i24.GSR = "ENABLED";
    FD1S3IX count_2170__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i25.GSR = "ENABLED";
    FD1S3IX count_2170__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i26.GSR = "ENABLED";
    FD1S3IX count_2170__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i27.GSR = "ENABLED";
    FD1S3IX count_2170__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i28.GSR = "ENABLED";
    FD1S3IX count_2170__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i29.GSR = "ENABLED";
    FD1S3IX count_2170__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i30.GSR = "ENABLED";
    FD1S3IX count_2170__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n28891), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2170__i31.GSR = "ENABLED";
    CCU2D sub_1722_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24041), .COUT(n24042));
    defparam sub_1722_add_2_3.INIT0 = 16'h5999;
    defparam sub_1722_add_2_3.INIT1 = 16'h5999;
    defparam sub_1722_add_2_3.INJECT1_0 = "NO";
    defparam sub_1722_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n24041));
    defparam sub_1722_add_2_1.INIT0 = 16'h0000;
    defparam sub_1722_add_2_1.INIT1 = 16'h5999;
    defparam sub_1722_add_2_1.INJECT1_0 = "NO";
    defparam sub_1722_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24040), .S1(n7086));
    defparam sub_1723_add_2_33.INIT0 = 16'hf555;
    defparam sub_1723_add_2_33.INIT1 = 16'h0000;
    defparam sub_1723_add_2_33.INJECT1_0 = "NO";
    defparam sub_1723_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24039), .COUT(n24040));
    defparam sub_1723_add_2_31.INIT0 = 16'hf555;
    defparam sub_1723_add_2_31.INIT1 = 16'hf555;
    defparam sub_1723_add_2_31.INJECT1_0 = "NO";
    defparam sub_1723_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24038), .COUT(n24039));
    defparam sub_1723_add_2_29.INIT0 = 16'hf555;
    defparam sub_1723_add_2_29.INIT1 = 16'hf555;
    defparam sub_1723_add_2_29.INJECT1_0 = "NO";
    defparam sub_1723_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24037), .COUT(n24038));
    defparam sub_1723_add_2_27.INIT0 = 16'hf555;
    defparam sub_1723_add_2_27.INIT1 = 16'hf555;
    defparam sub_1723_add_2_27.INJECT1_0 = "NO";
    defparam sub_1723_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24036), .COUT(n24037));
    defparam sub_1723_add_2_25.INIT0 = 16'hf555;
    defparam sub_1723_add_2_25.INIT1 = 16'hf555;
    defparam sub_1723_add_2_25.INJECT1_0 = "NO";
    defparam sub_1723_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24035), .COUT(n24036));
    defparam sub_1723_add_2_23.INIT0 = 16'hf555;
    defparam sub_1723_add_2_23.INIT1 = 16'hf555;
    defparam sub_1723_add_2_23.INJECT1_0 = "NO";
    defparam sub_1723_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24034), .COUT(n24035));
    defparam sub_1723_add_2_21.INIT0 = 16'hf555;
    defparam sub_1723_add_2_21.INIT1 = 16'hf555;
    defparam sub_1723_add_2_21.INJECT1_0 = "NO";
    defparam sub_1723_add_2_21.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n28891), .CD(n14373), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    CCU2D sub_1723_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24033), .COUT(n24034));
    defparam sub_1723_add_2_19.INIT0 = 16'hf555;
    defparam sub_1723_add_2_19.INIT1 = 16'hf555;
    defparam sub_1723_add_2_19.INJECT1_0 = "NO";
    defparam sub_1723_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24032), .COUT(n24033));
    defparam sub_1723_add_2_17.INIT0 = 16'hf555;
    defparam sub_1723_add_2_17.INIT1 = 16'hf555;
    defparam sub_1723_add_2_17.INJECT1_0 = "NO";
    defparam sub_1723_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24031), .COUT(n24032));
    defparam sub_1723_add_2_15.INIT0 = 16'hf555;
    defparam sub_1723_add_2_15.INIT1 = 16'hf555;
    defparam sub_1723_add_2_15.INJECT1_0 = "NO";
    defparam sub_1723_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24030), .COUT(n24031));
    defparam sub_1723_add_2_13.INIT0 = 16'hf555;
    defparam sub_1723_add_2_13.INIT1 = 16'hf555;
    defparam sub_1723_add_2_13.INJECT1_0 = "NO";
    defparam sub_1723_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24029), .COUT(n24030));
    defparam sub_1723_add_2_11.INIT0 = 16'hf555;
    defparam sub_1723_add_2_11.INIT1 = 16'hf555;
    defparam sub_1723_add_2_11.INJECT1_0 = "NO";
    defparam sub_1723_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24028), .COUT(n24029));
    defparam sub_1723_add_2_9.INIT0 = 16'hf555;
    defparam sub_1723_add_2_9.INIT1 = 16'hf555;
    defparam sub_1723_add_2_9.INJECT1_0 = "NO";
    defparam sub_1723_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24027), .COUT(n24028));
    defparam sub_1723_add_2_7.INIT0 = 16'hf555;
    defparam sub_1723_add_2_7.INIT1 = 16'hf555;
    defparam sub_1723_add_2_7.INJECT1_0 = "NO";
    defparam sub_1723_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24026), .COUT(n24027));
    defparam sub_1723_add_2_5.INIT0 = 16'hf555;
    defparam sub_1723_add_2_5.INIT1 = 16'hf555;
    defparam sub_1723_add_2_5.INJECT1_0 = "NO";
    defparam sub_1723_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24025), .COUT(n24026));
    defparam sub_1723_add_2_3.INIT0 = 16'hf555;
    defparam sub_1723_add_2_3.INIT1 = 16'hf555;
    defparam sub_1723_add_2_3.INJECT1_0 = "NO";
    defparam sub_1723_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1723_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n24025));
    defparam sub_1723_add_2_1.INIT0 = 16'h0000;
    defparam sub_1723_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1723_add_2_1.INJECT1_0 = "NO";
    defparam sub_1723_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1720_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24072), .S1(n7017));
    defparam sub_1720_add_2_33.INIT0 = 16'h5555;
    defparam sub_1720_add_2_33.INIT1 = 16'h0000;
    defparam sub_1720_add_2_33.INJECT1_0 = "NO";
    defparam sub_1720_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1720_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24071), .COUT(n24072));
    defparam sub_1720_add_2_31.INIT0 = 16'h5999;
    defparam sub_1720_add_2_31.INIT1 = 16'h5999;
    defparam sub_1720_add_2_31.INJECT1_0 = "NO";
    defparam sub_1720_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1720_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24070), .COUT(n24071));
    defparam sub_1720_add_2_29.INIT0 = 16'h5999;
    defparam sub_1720_add_2_29.INIT1 = 16'h5999;
    defparam sub_1720_add_2_29.INJECT1_0 = "NO";
    defparam sub_1720_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1720_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24069), .COUT(n24070));
    defparam sub_1720_add_2_27.INIT0 = 16'h5999;
    defparam sub_1720_add_2_27.INIT1 = 16'h5999;
    defparam sub_1720_add_2_27.INJECT1_0 = "NO";
    defparam sub_1720_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1720_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24068), .COUT(n24069));
    defparam sub_1720_add_2_25.INIT0 = 16'h5999;
    defparam sub_1720_add_2_25.INIT1 = 16'h5999;
    defparam sub_1720_add_2_25.INJECT1_0 = "NO";
    defparam sub_1720_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1720_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24067), .COUT(n24068));
    defparam sub_1720_add_2_23.INIT0 = 16'h5999;
    defparam sub_1720_add_2_23.INIT1 = 16'h5999;
    defparam sub_1720_add_2_23.INJECT1_0 = "NO";
    defparam sub_1720_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1720_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24066), .COUT(n24067));
    defparam sub_1720_add_2_21.INIT0 = 16'h5999;
    defparam sub_1720_add_2_21.INIT1 = 16'h5999;
    defparam sub_1720_add_2_21.INJECT1_0 = "NO";
    defparam sub_1720_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1720_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24065), .COUT(n24066));
    defparam sub_1720_add_2_19.INIT0 = 16'h5999;
    defparam sub_1720_add_2_19.INIT1 = 16'h5999;
    defparam sub_1720_add_2_19.INJECT1_0 = "NO";
    defparam sub_1720_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1720_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24064), .COUT(n24065));
    defparam sub_1720_add_2_17.INIT0 = 16'h5999;
    defparam sub_1720_add_2_17.INIT1 = 16'h5999;
    defparam sub_1720_add_2_17.INJECT1_0 = "NO";
    defparam sub_1720_add_2_17.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module ClockDivider_U10
//

module ClockDivider_U10 (debug_c_c, n241, n30647, n6670, n27582, n24993, 
            n28893, n27493, n24976, GND_net, n27569, n24988, n27575, 
            n24998, n27590, n24991, n27548, n11996, n27556, n11997, 
            n1018, n6, n27509, n26690, n27527, n12104, n27640, 
            n12804, n27638, n12807) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n241;
    input n30647;
    output n6670;
    input n27582;
    output n24993;
    output n28893;
    input n27493;
    output n24976;
    input GND_net;
    input n27569;
    output n24988;
    input n27575;
    output n24998;
    input n27590;
    output n24991;
    input n27548;
    output n11996;
    input n27556;
    output n11997;
    input n1018;
    output n6;
    input n27509;
    output n26690;
    input n27527;
    output n12104;
    input n27640;
    output n12804;
    input n27638;
    output n12807;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire clk_255kHz, n6705, n2546;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n24475, n24474, n24473, n24472, n24471, n24470, n24469, 
        n24468, n24467, n24466, n24465, n24216, n24464, n24463, 
        n24215, n24462, n24214, n24213, n24461, n24460, n24212, 
        n24211, n24210, n24209, n24208, n24207, n24206, n24205, 
        n24204, n24203, n24202, n24201, n24435, n24434, n24433, 
        n24432, n24431, n24430, n24429, n24428, n24427, n24426, 
        n24425, n24424, n24423, n24422, n24421;
    
    FD1S3AX clk_o_22 (.D(n241), .CK(debug_c_c), .Q(clk_255kHz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=508, LSE_RLINE=511 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    LUT4 i21300_2_lut_4_lut (.A(n30647), .B(clk_255kHz), .C(n6670), .D(n27582), 
         .Z(n24993)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21300_2_lut_4_lut.init = 16'h1000;
    LUT4 i889_2_lut (.A(n6705), .B(n30647), .Z(n2546)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i889_2_lut.init = 16'heeee;
    FD1S3IX count_2166__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2546), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i0.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_235 (.A(n30647), .B(clk_255kHz), .C(n6670), .Z(n28893)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i2_3_lut_rep_235.init = 16'h1010;
    LUT4 i21211_2_lut_4_lut (.A(n30647), .B(clk_255kHz), .C(n6670), .D(n27493), 
         .Z(n24976)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21211_2_lut_4_lut.init = 16'h1000;
    CCU2D count_2166_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24475), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_33.INIT1 = 16'h0000;
    defparam count_2166_add_4_33.INJECT1_0 = "NO";
    defparam count_2166_add_4_33.INJECT1_1 = "NO";
    LUT4 i21287_2_lut_4_lut (.A(n30647), .B(clk_255kHz), .C(n6670), .D(n27569), 
         .Z(n24988)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21287_2_lut_4_lut.init = 16'h1000;
    LUT4 i21293_2_lut_4_lut (.A(n30647), .B(clk_255kHz), .C(n6670), .D(n27575), 
         .Z(n24998)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21293_2_lut_4_lut.init = 16'h1000;
    CCU2D count_2166_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24474), .COUT(n24475), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2166_add_4_31.INJECT1_0 = "NO";
    defparam count_2166_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2166_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24473), .COUT(n24474), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2166_add_4_29.INJECT1_0 = "NO";
    defparam count_2166_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2166_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24472), .COUT(n24473), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2166_add_4_27.INJECT1_0 = "NO";
    defparam count_2166_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2166_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24471), .COUT(n24472), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2166_add_4_25.INJECT1_0 = "NO";
    defparam count_2166_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2166_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24470), .COUT(n24471), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2166_add_4_23.INJECT1_0 = "NO";
    defparam count_2166_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2166_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24469), .COUT(n24470), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2166_add_4_21.INJECT1_0 = "NO";
    defparam count_2166_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2166_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24468), .COUT(n24469), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2166_add_4_19.INJECT1_0 = "NO";
    defparam count_2166_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2166_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24467), .COUT(n24468), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2166_add_4_17.INJECT1_0 = "NO";
    defparam count_2166_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2166_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24466), .COUT(n24467), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2166_add_4_15.INJECT1_0 = "NO";
    defparam count_2166_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2166_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24465), .COUT(n24466), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2166_add_4_13.INJECT1_0 = "NO";
    defparam count_2166_add_4_13.INJECT1_1 = "NO";
    CCU2D sub_1705_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24216), .S0(n6705));
    defparam sub_1705_add_2_cout.INIT0 = 16'h0000;
    defparam sub_1705_add_2_cout.INIT1 = 16'h0000;
    defparam sub_1705_add_2_cout.INJECT1_0 = "NO";
    defparam sub_1705_add_2_cout.INJECT1_1 = "NO";
    CCU2D count_2166_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24464), .COUT(n24465), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2166_add_4_11.INJECT1_0 = "NO";
    defparam count_2166_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2166_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24463), .COUT(n24464), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2166_add_4_9.INJECT1_0 = "NO";
    defparam count_2166_add_4_9.INJECT1_1 = "NO";
    CCU2D sub_1705_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24215), .COUT(n24216));
    defparam sub_1705_add_2_32.INIT0 = 16'h5555;
    defparam sub_1705_add_2_32.INIT1 = 16'h5555;
    defparam sub_1705_add_2_32.INJECT1_0 = "NO";
    defparam sub_1705_add_2_32.INJECT1_1 = "NO";
    CCU2D count_2166_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24462), .COUT(n24463), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2166_add_4_7.INJECT1_0 = "NO";
    defparam count_2166_add_4_7.INJECT1_1 = "NO";
    CCU2D sub_1705_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24214), .COUT(n24215));
    defparam sub_1705_add_2_30.INIT0 = 16'h5555;
    defparam sub_1705_add_2_30.INIT1 = 16'h5555;
    defparam sub_1705_add_2_30.INJECT1_0 = "NO";
    defparam sub_1705_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_1705_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24213), .COUT(n24214));
    defparam sub_1705_add_2_28.INIT0 = 16'h5555;
    defparam sub_1705_add_2_28.INIT1 = 16'h5555;
    defparam sub_1705_add_2_28.INJECT1_0 = "NO";
    defparam sub_1705_add_2_28.INJECT1_1 = "NO";
    LUT4 i21308_2_lut_4_lut (.A(n30647), .B(clk_255kHz), .C(n6670), .D(n27590), 
         .Z(n24991)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21308_2_lut_4_lut.init = 16'h1000;
    CCU2D count_2166_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24461), .COUT(n24462), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2166_add_4_5.INJECT1_0 = "NO";
    defparam count_2166_add_4_5.INJECT1_1 = "NO";
    LUT4 i21266_2_lut_4_lut (.A(n30647), .B(clk_255kHz), .C(n6670), .D(n27548), 
         .Z(n11996)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21266_2_lut_4_lut.init = 16'h1000;
    LUT4 i21274_2_lut_4_lut (.A(n30647), .B(clk_255kHz), .C(n6670), .D(n27556), 
         .Z(n11997)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21274_2_lut_4_lut.init = 16'h1000;
    CCU2D count_2166_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24460), .COUT(n24461), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2166_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2166_add_4_3.INJECT1_0 = "NO";
    defparam count_2166_add_4_3.INJECT1_1 = "NO";
    LUT4 i2_2_lut_4_lut (.A(n30647), .B(clk_255kHz), .C(n6670), .D(n1018), 
         .Z(n6)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i2_2_lut_4_lut.init = 16'h1000;
    LUT4 i21227_2_lut_4_lut (.A(n30647), .B(clk_255kHz), .C(n6670), .D(n27509), 
         .Z(n26690)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21227_2_lut_4_lut.init = 16'h1000;
    CCU2D count_2166_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24460), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166_add_4_1.INIT0 = 16'hF000;
    defparam count_2166_add_4_1.INIT1 = 16'h0555;
    defparam count_2166_add_4_1.INJECT1_0 = "NO";
    defparam count_2166_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_1705_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24212), .COUT(n24213));
    defparam sub_1705_add_2_26.INIT0 = 16'h5555;
    defparam sub_1705_add_2_26.INIT1 = 16'h5555;
    defparam sub_1705_add_2_26.INJECT1_0 = "NO";
    defparam sub_1705_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_1705_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24211), .COUT(n24212));
    defparam sub_1705_add_2_24.INIT0 = 16'h5555;
    defparam sub_1705_add_2_24.INIT1 = 16'h5555;
    defparam sub_1705_add_2_24.INJECT1_0 = "NO";
    defparam sub_1705_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_1705_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24210), .COUT(n24211));
    defparam sub_1705_add_2_22.INIT0 = 16'h5555;
    defparam sub_1705_add_2_22.INIT1 = 16'h5555;
    defparam sub_1705_add_2_22.INJECT1_0 = "NO";
    defparam sub_1705_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_1705_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24209), .COUT(n24210));
    defparam sub_1705_add_2_20.INIT0 = 16'h5555;
    defparam sub_1705_add_2_20.INIT1 = 16'h5555;
    defparam sub_1705_add_2_20.INJECT1_0 = "NO";
    defparam sub_1705_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_1705_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24208), .COUT(n24209));
    defparam sub_1705_add_2_18.INIT0 = 16'h5555;
    defparam sub_1705_add_2_18.INIT1 = 16'h5555;
    defparam sub_1705_add_2_18.INJECT1_0 = "NO";
    defparam sub_1705_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_1705_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24207), .COUT(n24208));
    defparam sub_1705_add_2_16.INIT0 = 16'h5555;
    defparam sub_1705_add_2_16.INIT1 = 16'h5555;
    defparam sub_1705_add_2_16.INJECT1_0 = "NO";
    defparam sub_1705_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_1705_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24206), .COUT(n24207));
    defparam sub_1705_add_2_14.INIT0 = 16'h5555;
    defparam sub_1705_add_2_14.INIT1 = 16'h5555;
    defparam sub_1705_add_2_14.INJECT1_0 = "NO";
    defparam sub_1705_add_2_14.INJECT1_1 = "NO";
    LUT4 i21245_2_lut_4_lut (.A(n30647), .B(clk_255kHz), .C(n6670), .D(n27527), 
         .Z(n12104)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21245_2_lut_4_lut.init = 16'h1000;
    CCU2D sub_1705_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24205), .COUT(n24206));
    defparam sub_1705_add_2_12.INIT0 = 16'h5555;
    defparam sub_1705_add_2_12.INIT1 = 16'h5555;
    defparam sub_1705_add_2_12.INJECT1_0 = "NO";
    defparam sub_1705_add_2_12.INJECT1_1 = "NO";
    LUT4 i21358_2_lut_4_lut (.A(n30647), .B(clk_255kHz), .C(n6670), .D(n27640), 
         .Z(n12804)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21358_2_lut_4_lut.init = 16'h1000;
    CCU2D sub_1705_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24204), .COUT(n24205));
    defparam sub_1705_add_2_10.INIT0 = 16'h5555;
    defparam sub_1705_add_2_10.INIT1 = 16'h5555;
    defparam sub_1705_add_2_10.INJECT1_0 = "NO";
    defparam sub_1705_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_1705_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24203), .COUT(n24204));
    defparam sub_1705_add_2_8.INIT0 = 16'h5555;
    defparam sub_1705_add_2_8.INIT1 = 16'h5555;
    defparam sub_1705_add_2_8.INJECT1_0 = "NO";
    defparam sub_1705_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_1705_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24202), .COUT(n24203));
    defparam sub_1705_add_2_6.INIT0 = 16'h5555;
    defparam sub_1705_add_2_6.INIT1 = 16'h5aaa;
    defparam sub_1705_add_2_6.INJECT1_0 = "NO";
    defparam sub_1705_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_1705_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24201), .COUT(n24202));
    defparam sub_1705_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_1705_add_2_4.INIT1 = 16'h5aaa;
    defparam sub_1705_add_2_4.INJECT1_0 = "NO";
    defparam sub_1705_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_1705_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24201));
    defparam sub_1705_add_2_2.INIT0 = 16'h0000;
    defparam sub_1705_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_1705_add_2_2.INJECT1_0 = "NO";
    defparam sub_1705_add_2_2.INJECT1_1 = "NO";
    LUT4 i21356_2_lut_4_lut (.A(n30647), .B(clk_255kHz), .C(n6670), .D(n27638), 
         .Z(n12807)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i21356_2_lut_4_lut.init = 16'h1000;
    CCU2D add_18237_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24435), 
          .S1(n6670));
    defparam add_18237_32.INIT0 = 16'h5555;
    defparam add_18237_32.INIT1 = 16'h0000;
    defparam add_18237_32.INJECT1_0 = "NO";
    defparam add_18237_32.INJECT1_1 = "NO";
    FD1S3IX count_2166__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2546), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i1.GSR = "ENABLED";
    CCU2D add_18237_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24434), .COUT(n24435));
    defparam add_18237_30.INIT0 = 16'h5555;
    defparam add_18237_30.INIT1 = 16'h5555;
    defparam add_18237_30.INJECT1_0 = "NO";
    defparam add_18237_30.INJECT1_1 = "NO";
    CCU2D add_18237_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24433), .COUT(n24434));
    defparam add_18237_28.INIT0 = 16'h5555;
    defparam add_18237_28.INIT1 = 16'h5555;
    defparam add_18237_28.INJECT1_0 = "NO";
    defparam add_18237_28.INJECT1_1 = "NO";
    FD1S3IX count_2166__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2546), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i2.GSR = "ENABLED";
    FD1S3IX count_2166__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2546), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i3.GSR = "ENABLED";
    FD1S3IX count_2166__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2546), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i4.GSR = "ENABLED";
    FD1S3IX count_2166__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2546), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i5.GSR = "ENABLED";
    FD1S3IX count_2166__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2546), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i6.GSR = "ENABLED";
    FD1S3IX count_2166__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2546), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i7.GSR = "ENABLED";
    FD1S3IX count_2166__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2546), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i8.GSR = "ENABLED";
    FD1S3IX count_2166__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2546), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i9.GSR = "ENABLED";
    FD1S3IX count_2166__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i10.GSR = "ENABLED";
    FD1S3IX count_2166__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i11.GSR = "ENABLED";
    FD1S3IX count_2166__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i12.GSR = "ENABLED";
    FD1S3IX count_2166__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i13.GSR = "ENABLED";
    FD1S3IX count_2166__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i14.GSR = "ENABLED";
    FD1S3IX count_2166__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i15.GSR = "ENABLED";
    FD1S3IX count_2166__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i16.GSR = "ENABLED";
    FD1S3IX count_2166__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i17.GSR = "ENABLED";
    FD1S3IX count_2166__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i18.GSR = "ENABLED";
    FD1S3IX count_2166__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i19.GSR = "ENABLED";
    FD1S3IX count_2166__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i20.GSR = "ENABLED";
    FD1S3IX count_2166__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i21.GSR = "ENABLED";
    FD1S3IX count_2166__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i22.GSR = "ENABLED";
    FD1S3IX count_2166__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i23.GSR = "ENABLED";
    FD1S3IX count_2166__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i24.GSR = "ENABLED";
    FD1S3IX count_2166__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i25.GSR = "ENABLED";
    FD1S3IX count_2166__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i26.GSR = "ENABLED";
    FD1S3IX count_2166__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i27.GSR = "ENABLED";
    FD1S3IX count_2166__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i28.GSR = "ENABLED";
    FD1S3IX count_2166__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i29.GSR = "ENABLED";
    FD1S3IX count_2166__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i30.GSR = "ENABLED";
    FD1S3IX count_2166__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2546), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2166__i31.GSR = "ENABLED";
    CCU2D add_18237_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24432), .COUT(n24433));
    defparam add_18237_26.INIT0 = 16'h5555;
    defparam add_18237_26.INIT1 = 16'h5555;
    defparam add_18237_26.INJECT1_0 = "NO";
    defparam add_18237_26.INJECT1_1 = "NO";
    CCU2D add_18237_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24431), .COUT(n24432));
    defparam add_18237_24.INIT0 = 16'h5555;
    defparam add_18237_24.INIT1 = 16'h5555;
    defparam add_18237_24.INJECT1_0 = "NO";
    defparam add_18237_24.INJECT1_1 = "NO";
    CCU2D add_18237_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24430), .COUT(n24431));
    defparam add_18237_22.INIT0 = 16'h5555;
    defparam add_18237_22.INIT1 = 16'h5555;
    defparam add_18237_22.INJECT1_0 = "NO";
    defparam add_18237_22.INJECT1_1 = "NO";
    CCU2D add_18237_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24429), .COUT(n24430));
    defparam add_18237_20.INIT0 = 16'h5555;
    defparam add_18237_20.INIT1 = 16'h5555;
    defparam add_18237_20.INJECT1_0 = "NO";
    defparam add_18237_20.INJECT1_1 = "NO";
    CCU2D add_18237_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24428), .COUT(n24429));
    defparam add_18237_18.INIT0 = 16'h5555;
    defparam add_18237_18.INIT1 = 16'h5555;
    defparam add_18237_18.INJECT1_0 = "NO";
    defparam add_18237_18.INJECT1_1 = "NO";
    CCU2D add_18237_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24427), .COUT(n24428));
    defparam add_18237_16.INIT0 = 16'h5555;
    defparam add_18237_16.INIT1 = 16'h5555;
    defparam add_18237_16.INJECT1_0 = "NO";
    defparam add_18237_16.INJECT1_1 = "NO";
    CCU2D add_18237_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24426), .COUT(n24427));
    defparam add_18237_14.INIT0 = 16'h5555;
    defparam add_18237_14.INIT1 = 16'h5555;
    defparam add_18237_14.INJECT1_0 = "NO";
    defparam add_18237_14.INJECT1_1 = "NO";
    CCU2D add_18237_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24425), .COUT(n24426));
    defparam add_18237_12.INIT0 = 16'h5555;
    defparam add_18237_12.INIT1 = 16'h5555;
    defparam add_18237_12.INJECT1_0 = "NO";
    defparam add_18237_12.INJECT1_1 = "NO";
    CCU2D add_18237_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24424), .COUT(n24425));
    defparam add_18237_10.INIT0 = 16'h5555;
    defparam add_18237_10.INIT1 = 16'h5555;
    defparam add_18237_10.INJECT1_0 = "NO";
    defparam add_18237_10.INJECT1_1 = "NO";
    CCU2D add_18237_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24423), 
          .COUT(n24424));
    defparam add_18237_8.INIT0 = 16'h5555;
    defparam add_18237_8.INIT1 = 16'h5555;
    defparam add_18237_8.INJECT1_0 = "NO";
    defparam add_18237_8.INJECT1_1 = "NO";
    CCU2D add_18237_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24422), 
          .COUT(n24423));
    defparam add_18237_6.INIT0 = 16'h5555;
    defparam add_18237_6.INIT1 = 16'h5555;
    defparam add_18237_6.INJECT1_0 = "NO";
    defparam add_18237_6.INJECT1_1 = "NO";
    CCU2D add_18237_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24421), 
          .COUT(n24422));
    defparam add_18237_4.INIT0 = 16'h5555;
    defparam add_18237_4.INIT1 = 16'h5aaa;
    defparam add_18237_4.INJECT1_0 = "NO";
    defparam add_18237_4.INJECT1_1 = "NO";
    CCU2D add_18237_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24421));
    defparam add_18237_2.INIT0 = 16'h7000;
    defparam add_18237_2.INIT1 = 16'h5aaa;
    defparam add_18237_2.INJECT1_0 = "NO";
    defparam add_18237_2.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0) 
//

module \ArmPeripheral(axis_haddr=8'b0)  (\register_addr[1] , \register_addr[0] , 
            databus, n3446, read_value, debug_c_c, n11908, GND_net, 
            n30651, n30648, n30649, \read_size[0] , n28920, Stepper_X_M0_c_0, 
            n580, prev_select, n28927, n30650, \steps_reg[7] , n30652, 
            n609, n611, \control_reg[7] , n574, Stepper_X_Dir_c, Stepper_X_M2_c_2, 
            Stepper_X_M1_c_1, \read_size[2] , n28901, n30653, n28991, 
            rw, n28903, n29052, n28917, Stepper_X_En_c, Stepper_X_Step_c, 
            limit_c_0, n29025, n30647, n28898, n28965, n24994, n21, 
            VCC_net, Stepper_X_nFault_c, n13) /* synthesis syn_module_defined=1 */ ;
    input \register_addr[1] ;
    input \register_addr[0] ;
    input [31:0]databus;
    input n3446;
    output [31:0]read_value;
    input debug_c_c;
    input n11908;
    input GND_net;
    input n30651;
    input n30648;
    input n30649;
    output \read_size[0] ;
    input n28920;
    output Stepper_X_M0_c_0;
    input n580;
    output prev_select;
    input n28927;
    input n30650;
    output \steps_reg[7] ;
    input n30652;
    input n609;
    input n611;
    output \control_reg[7] ;
    input n574;
    output Stepper_X_Dir_c;
    output Stepper_X_M2_c_2;
    output Stepper_X_M1_c_1;
    output \read_size[2] ;
    input n28901;
    input n30653;
    input n28991;
    input rw;
    input n28903;
    input n29052;
    input n28917;
    output Stepper_X_En_c;
    output Stepper_X_Step_c;
    input limit_c_0;
    input n29025;
    input n30647;
    input n28898;
    input n28965;
    output n24994;
    input n21;
    input VCC_net;
    input Stepper_X_nFault_c;
    input n13;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire n26880;
    wire [31:0]n225;
    wire [31:0]n3447;
    wire [31:0]n5184;
    
    wire n26894, n12075, prev_step_clk, step_clk, limit_latched, n183, 
        prev_limit_latched, n12444, n1, n2, n1_adj_249, n2_adj_250, 
        n1_adj_251, n2_adj_252, n1_adj_253, n2_adj_254, int_step, 
        n12, n28908, n28896, n28897, n9604;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n17333, n27430, n26895, n27431, fault_latched, n27433, 
        n27434, n26885, n26884, n26883, n26882, n26881, n27439, 
        n27440, n27441, n49, n62, n58, n50, n41, n60, n54, 
        n42, n52, n38, n56, n46, n27432, n27435, n26879, n26878, 
        n24420, n24419, n24418, n26872, n26876, n26874, n26875, 
        n26873, n26877, n26887, n26886, n26888, n26889, n26890, 
        n26891, n24417, n26892, n26893, n24416, n24415, n24414, 
        n24413, n24412, n24411, n24410, n24409, n24408, n24407, 
        n24406, n24405;
    
    LUT4 i1_4_lut (.A(div_factor_reg[13]), .B(\register_addr[1] ), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n26880)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 mux_1380_i10_3_lut (.A(n225[9]), .B(databus[9]), .C(n3446), .Z(n3447[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i9_3_lut (.A(n225[8]), .B(databus[8]), .C(n3446), .Z(n3447[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i9_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i5 (.D(n5184[5]), .SP(n11908), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    LUT4 mux_1380_i8_3_lut (.A(n225[7]), .B(databus[7]), .C(n3446), .Z(n3447[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i8_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i19 (.D(n3447[19]), .CK(debug_c_c), .CD(n30651), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_165 (.A(div_factor_reg[30]), .B(\register_addr[1] ), 
         .C(steps_reg[30]), .D(\register_addr[0] ), .Z(n26894)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_165.init = 16'hc088;
    FD1S3IX steps_reg__i18 (.D(n3447[18]), .CK(debug_c_c), .CD(n30648), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3447[17]), .CK(debug_c_c), .CD(n30648), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3447[16]), .CK(debug_c_c), .CD(n30648), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3447[0]), .CK(debug_c_c), .CD(n30648), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3447[15]), .CK(debug_c_c), .CD(n30648), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3447[14]), .CK(debug_c_c), .CD(n30649), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n28920), .SP(n11908), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3447[13]), .CK(debug_c_c), .CD(n30649), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3447[12]), .CK(debug_c_c), .CD(n30649), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n580), .SP(n12075), .CK(debug_c_c), .Q(Stepper_X_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_176 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_176.GSR = "ENABLED";
    FD1S3AX limit_latched_177 (.D(n183), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_177.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_178 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_178.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n580), .SP(n12444), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3447[11]), .CK(debug_c_c), .CD(n30649), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3AX prev_select_175 (.D(n28927), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_175.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3447[10]), .CK(debug_c_c), .CD(n30649), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    LUT4 mux_1380_i7_3_lut (.A(n225[6]), .B(databus[6]), .C(n3446), .Z(n3447[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i7_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i9 (.D(n3447[9]), .CK(debug_c_c), .CD(n30649), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3447[8]), .CK(debug_c_c), .CD(n30650), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3447[7]), .CK(debug_c_c), .CD(n30650), 
            .Q(\steps_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3447[6]), .CK(debug_c_c), .CD(n30650), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    PFUMX mux_1596_Mux_3_i3 (.BLUT(n1), .ALUT(n2), .C0(\register_addr[1] ), 
          .Z(n5184[3]));
    PFUMX mux_1596_Mux_4_i3 (.BLUT(n1_adj_249), .ALUT(n2_adj_250), .C0(\register_addr[1] ), 
          .Z(n5184[4]));
    FD1S3IX steps_reg__i5 (.D(n3447[5]), .CK(debug_c_c), .CD(n30650), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3447[4]), .CK(debug_c_c), .CD(n30650), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3447[3]), .CK(debug_c_c), .CD(n30650), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3447[2]), .CK(debug_c_c), .CD(n30650), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3447[1]), .CK(debug_c_c), .CD(n30650), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    PFUMX mux_1596_Mux_5_i3 (.BLUT(n1_adj_251), .ALUT(n2_adj_252), .C0(\register_addr[1] ), 
          .Z(n5184[5]));
    PFUMX mux_1596_Mux_6_i3 (.BLUT(n1_adj_253), .ALUT(n2_adj_254), .C0(\register_addr[1] ), 
          .Z(n5184[6]));
    FD1P3AX int_step_183 (.D(n28908), .SP(n12), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_183.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n28896), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n28896), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n28896), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n28896), .PD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n28896), .PD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n28896), .PD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n28896), .PD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n28896), .PD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n28896), .PD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n28896), .PD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n609), .SP(n12444), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n611), .SP(n12444), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n28896), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n28897), .CD(n9604), .CK(debug_c_c), 
            .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3AX control_reg_i7 (.D(n574), .SP(n12075), .CK(debug_c_c), .Q(control_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n28897), .PD(n30652), 
            .CK(debug_c_c), .Q(Stepper_X_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n609), .SP(n12075), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n28897), .PD(n30652), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n611), .SP(n12075), .CK(debug_c_c), .Q(Stepper_X_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n28897), .PD(n30652), 
            .CK(debug_c_c), .Q(Stepper_X_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n28901), .SP(n11908), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3447[31]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3447[30]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3447[29]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3447[28]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3447[27]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3447[26]), .CK(debug_c_c), .CD(n30653), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3447[25]), .CK(debug_c_c), .CD(n28991), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3447[24]), .CK(debug_c_c), .CD(n28991), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3447[23]), .CK(debug_c_c), .CD(n28991), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3447[22]), .CK(debug_c_c), .CD(n28991), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3447[21]), .CK(debug_c_c), .CD(n28991), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3447[20]), .CK(debug_c_c), .CD(n28991), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n12444), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n12444), .CD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n12444), .CD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n12444), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n12444), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n12444), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n12444), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n12444), .CD(n30651), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n12444), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n12444), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n12444), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n12444), .CD(n30648), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n12444), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n12444), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n12444), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n12444), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n12444), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n12444), .CD(n30652), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    LUT4 i11582_3_lut (.A(\control_reg[7] ), .B(div_factor_reg[7]), .C(\register_addr[1] ), 
         .Z(n17333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i11582_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i18_3_lut (.A(n225[17]), .B(databus[17]), .C(n3446), 
         .Z(n3447[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i17_3_lut (.A(n225[16]), .B(databus[16]), .C(n3446), 
         .Z(n3447[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i17_3_lut.init = 16'hcaca;
    LUT4 i14314_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n1)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14314_2_lut.init = 16'h2222;
    LUT4 mux_1380_i1_3_lut (.A(n225[0]), .B(databus[0]), .C(n3446), .Z(n3447[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i1_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_238_4_lut (.A(rw), .B(n28903), .C(n29052), .D(n28917), 
         .Z(n28896)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i2_3_lut_rep_238_4_lut.init = 16'h0040;
    LUT4 mux_1380_i16_3_lut (.A(n225[15]), .B(databus[15]), .C(n3446), 
         .Z(n3447[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i15_3_lut (.A(n225[14]), .B(databus[14]), .C(n3446), 
         .Z(n3447[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1596_Mux_3_i2_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), 
         .C(\register_addr[0] ), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1596_Mux_3_i2_3_lut.init = 16'hcaca;
    LUT4 i14313_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n1_adj_249)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14313_2_lut.init = 16'h2222;
    LUT4 i11589_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n2_adj_250)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i11589_3_lut.init = 16'hcaca;
    LUT4 i8_1_lut (.A(control_reg[6]), .Z(Stepper_X_En_c)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(44[14:29])
    defparam i8_1_lut.init = 16'h5555;
    LUT4 i1_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_X_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 mux_1380_i6_3_lut (.A(n225[5]), .B(databus[5]), .C(n3446), .Z(n3447[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i5_3_lut (.A(n225[4]), .B(databus[4]), .C(n3446), .Z(n3447[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i4_3_lut (.A(n225[3]), .B(databus[3]), .C(n3446), .Z(n3447[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i14_3_lut (.A(n225[13]), .B(databus[13]), .C(n3446), 
         .Z(n3447[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i3_3_lut (.A(n225[2]), .B(databus[2]), .C(n3446), .Z(n3447[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i2_3_lut (.A(n225[1]), .B(databus[1]), .C(n3446), .Z(n3447[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i2_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i6 (.D(n5184[6]), .SP(n11908), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    LUT4 mux_1380_i13_3_lut (.A(n225[12]), .B(databus[12]), .C(n3446), 
         .Z(n3447[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i13_3_lut.init = 16'hcaca;
    LUT4 i14312_2_lut (.A(Stepper_X_Dir_c), .B(\register_addr[0] ), .Z(n1_adj_251)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14312_2_lut.init = 16'h2222;
    LUT4 mux_1596_Mux_5_i2_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), 
         .C(\register_addr[0] ), .Z(n2_adj_252)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1596_Mux_5_i2_3_lut.init = 16'hcaca;
    LUT4 i14311_2_lut (.A(control_reg[6]), .B(\register_addr[0] ), .Z(n1_adj_253)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14311_2_lut.init = 16'h2222;
    LUT4 i21060_3_lut (.A(Stepper_X_M2_c_2), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n27430)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21060_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_166 (.A(div_factor_reg[31]), .B(\register_addr[1] ), 
         .C(steps_reg[31]), .D(\register_addr[0] ), .Z(n26895)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_166.init = 16'hc088;
    LUT4 mux_1596_Mux_6_i2_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), 
         .C(\register_addr[0] ), .Z(n2_adj_254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1596_Mux_6_i2_3_lut.init = 16'hcaca;
    LUT4 i21061_3_lut (.A(div_factor_reg[2]), .B(steps_reg[2]), .C(\register_addr[0] ), 
         .Z(n27431)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21061_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i7 (.D(n5184[7]), .SP(n11908), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    LUT4 i21063_3_lut (.A(Stepper_X_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n27433)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21063_3_lut.init = 16'hcaca;
    LUT4 i21064_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n27434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21064_3_lut.init = 16'hcaca;
    LUT4 i119_1_lut (.A(limit_c_0), .Z(n183)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i119_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_167 (.A(div_factor_reg[8]), .B(\register_addr[1] ), 
         .C(steps_reg[8]), .D(\register_addr[0] ), .Z(n26885)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_167.init = 16'hc088;
    FD1P3AX read_value__i8 (.D(n26885), .SP(n11908), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    LUT4 mux_1380_i12_3_lut (.A(n225[11]), .B(databus[11]), .C(n3446), 
         .Z(n3447[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i11_3_lut (.A(n225[10]), .B(databus[10]), .C(n3446), 
         .Z(n3447[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i11_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i9 (.D(n26884), .SP(n11908), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n26883), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n26882), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n26881), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    PFUMX i21071 (.BLUT(n27439), .ALUT(n27440), .C0(\register_addr[0] ), 
          .Z(n27441));
    LUT4 i1_4_lut_adj_168 (.A(div_factor_reg[9]), .B(\register_addr[1] ), 
         .C(steps_reg[9]), .D(\register_addr[0] ), .Z(n26884)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_168.init = 16'hc088;
    LUT4 i1_4_lut_adj_169 (.A(div_factor_reg[10]), .B(\register_addr[1] ), 
         .C(steps_reg[10]), .D(\register_addr[0] ), .Z(n26883)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_169.init = 16'hc088;
    LUT4 i1_4_lut_adj_170 (.A(div_factor_reg[11]), .B(\register_addr[1] ), 
         .C(steps_reg[11]), .D(\register_addr[0] ), .Z(n26882)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_170.init = 16'hc088;
    FD1P3AX read_value__i13 (.D(n26880), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_171 (.A(div_factor_reg[12]), .B(\register_addr[1] ), 
         .C(steps_reg[12]), .D(\register_addr[0] ), .Z(n26881)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_171.init = 16'hc088;
    LUT4 i21360_2_lut_4_lut_4_lut (.A(n29025), .B(n30647), .C(n28898), 
         .D(n28965), .Z(n12075)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i21360_2_lut_4_lut_4_lut.init = 16'hccdc;
    LUT4 i21264_3_lut_rep_239_4_lut_4_lut (.A(n29025), .B(n28965), .C(n28903), 
         .D(rw), .Z(n28897)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i21264_3_lut_rep_239_4_lut_4_lut.init = 16'h0010;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n24994)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[8]), .B(steps_reg[18]), .C(steps_reg[28]), 
         .D(steps_reg[24]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[26]), .B(n52), .C(n38), .D(steps_reg[9]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[4]), .B(steps_reg[21]), .C(steps_reg[11]), 
         .D(steps_reg[25]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[30]), .B(\steps_reg[7] ), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[0]), .B(n56), .C(n46), .D(steps_reg[1]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[22]), .B(steps_reg[6]), .C(steps_reg[5]), 
         .D(steps_reg[10]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[14]), .B(steps_reg[19]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[29]), .B(steps_reg[3]), .C(steps_reg[13]), 
         .D(steps_reg[31]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[15]), .B(steps_reg[23]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[20]), .C(steps_reg[2]), 
         .D(steps_reg[27]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i21069_3_lut (.A(Stepper_X_M0_c_0), .B(div_factor_reg[0]), .C(\register_addr[1] ), 
         .Z(n27439)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21069_3_lut.init = 16'hcaca;
    PFUMX i21062 (.BLUT(n27430), .ALUT(n27431), .C0(\register_addr[1] ), 
          .Z(n27432));
    LUT4 i21070_3_lut (.A(n21), .B(steps_reg[0]), .C(\register_addr[1] ), 
         .Z(n27440)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21070_3_lut.init = 16'hcaca;
    PFUMX i21065 (.BLUT(n27433), .ALUT(n27434), .C0(\register_addr[1] ), 
          .Z(n27435));
    LUT4 mux_1380_i32_3_lut (.A(n225[31]), .B(databus[31]), .C(n3446), 
         .Z(n3447[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i32_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i0 (.D(n27441), .SP(n11908), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 mux_1380_i31_3_lut (.A(n225[30]), .B(databus[30]), .C(n3446), 
         .Z(n3447[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i30_3_lut (.A(n225[29]), .B(databus[29]), .C(n3446), 
         .Z(n3447[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i29_3_lut (.A(n225[28]), .B(databus[28]), .C(n3446), 
         .Z(n3447[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i28_3_lut (.A(n225[27]), .B(databus[27]), .C(n3446), 
         .Z(n3447[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i27_3_lut (.A(n225[26]), .B(databus[26]), .C(n3446), 
         .Z(n3447[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i19_3_lut (.A(n225[18]), .B(databus[18]), .C(n3446), 
         .Z(n3447[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i19_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i14 (.D(n26879), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n26878), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    IFS1P3DX fault_latched_179 (.D(Stepper_X_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_179.GSR = "ENABLED";
    CCU2D sub_126_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24420), .S0(n225[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_33.INIT0 = 16'h5555;
    defparam sub_126_add_2_33.INIT1 = 16'h0000;
    defparam sub_126_add_2_33.INJECT1_0 = "NO";
    defparam sub_126_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24419), .COUT(n24420), .S0(n225[29]), 
          .S1(n225[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_31.INIT0 = 16'h5555;
    defparam sub_126_add_2_31.INIT1 = 16'h5555;
    defparam sub_126_add_2_31.INJECT1_0 = "NO";
    defparam sub_126_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24418), .COUT(n24419), .S0(n225[27]), 
          .S1(n225[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_29.INIT0 = 16'h5555;
    defparam sub_126_add_2_29.INIT1 = 16'h5555;
    defparam sub_126_add_2_29.INJECT1_0 = "NO";
    defparam sub_126_add_2_29.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_172 (.A(div_factor_reg[14]), .B(\register_addr[1] ), 
         .C(steps_reg[14]), .D(\register_addr[0] ), .Z(n26879)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_172.init = 16'hc088;
    LUT4 i1_4_lut_adj_173 (.A(div_factor_reg[15]), .B(\register_addr[1] ), 
         .C(steps_reg[15]), .D(\register_addr[0] ), .Z(n26878)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_173.init = 16'hc088;
    FD1P3AX read_value__i16 (.D(n26872), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n26876), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n26874), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n26875), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n26873), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n26877), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n26887), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n26886), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n26888), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n26889), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n26890), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n26891), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    CCU2D sub_126_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24417), .COUT(n24418), .S0(n225[25]), 
          .S1(n225[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_27.INIT0 = 16'h5555;
    defparam sub_126_add_2_27.INIT1 = 16'h5555;
    defparam sub_126_add_2_27.INJECT1_0 = "NO";
    defparam sub_126_add_2_27.INJECT1_1 = "NO";
    FD1P3AX read_value__i28 (.D(n26892), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n26893), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n26894), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n26895), .SP(n11908), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    CCU2D sub_126_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24416), .COUT(n24417), .S0(n225[23]), 
          .S1(n225[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_25.INIT0 = 16'h5555;
    defparam sub_126_add_2_25.INIT1 = 16'h5555;
    defparam sub_126_add_2_25.INJECT1_0 = "NO";
    defparam sub_126_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24415), .COUT(n24416), .S0(n225[21]), 
          .S1(n225[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_23.INIT0 = 16'h5555;
    defparam sub_126_add_2_23.INIT1 = 16'h5555;
    defparam sub_126_add_2_23.INJECT1_0 = "NO";
    defparam sub_126_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24414), .COUT(n24415), .S0(n225[19]), 
          .S1(n225[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_21.INIT0 = 16'h5555;
    defparam sub_126_add_2_21.INIT1 = 16'h5555;
    defparam sub_126_add_2_21.INJECT1_0 = "NO";
    defparam sub_126_add_2_21.INJECT1_1 = "NO";
    LUT4 mux_1380_i26_3_lut (.A(n225[25]), .B(databus[25]), .C(n3446), 
         .Z(n3447[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i26_3_lut.init = 16'hcaca;
    CCU2D sub_126_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24413), .COUT(n24414), .S0(n225[17]), 
          .S1(n225[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_19.INIT0 = 16'h5555;
    defparam sub_126_add_2_19.INIT1 = 16'h5555;
    defparam sub_126_add_2_19.INJECT1_0 = "NO";
    defparam sub_126_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24412), .COUT(n24413), .S0(n225[15]), 
          .S1(n225[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_17.INIT0 = 16'h5555;
    defparam sub_126_add_2_17.INIT1 = 16'h5555;
    defparam sub_126_add_2_17.INJECT1_0 = "NO";
    defparam sub_126_add_2_17.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_174 (.A(div_factor_reg[16]), .B(\register_addr[1] ), 
         .C(steps_reg[16]), .D(\register_addr[0] ), .Z(n26872)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_174.init = 16'hc088;
    LUT4 mux_1380_i25_3_lut (.A(n225[24]), .B(databus[24]), .C(n3446), 
         .Z(n3447[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1380_i20_3_lut (.A(n225[19]), .B(databus[19]), .C(n3446), 
         .Z(n3447[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i20_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_175 (.A(div_factor_reg[17]), .B(\register_addr[1] ), 
         .C(steps_reg[17]), .D(\register_addr[0] ), .Z(n26876)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_175.init = 16'hc088;
    LUT4 i1_4_lut_adj_176 (.A(div_factor_reg[18]), .B(\register_addr[1] ), 
         .C(steps_reg[18]), .D(\register_addr[0] ), .Z(n26874)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_176.init = 16'hc088;
    FD1P3IX read_value__i1 (.D(n27435), .SP(n11908), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 mux_1380_i24_3_lut (.A(n225[23]), .B(databus[23]), .C(n3446), 
         .Z(n3447[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i24_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i2 (.D(n27432), .SP(n11908), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n5184[3]), .SP(n11908), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    LUT4 mux_1380_i23_3_lut (.A(n225[22]), .B(databus[22]), .C(n3446), 
         .Z(n3447[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i23_3_lut.init = 16'hcaca;
    PFUMX i11584 (.BLUT(n17333), .ALUT(n13), .C0(\register_addr[0] ), 
          .Z(n5184[7]));
    LUT4 i1_4_lut_adj_177 (.A(div_factor_reg[19]), .B(\register_addr[1] ), 
         .C(steps_reg[19]), .D(\register_addr[0] ), .Z(n26875)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_177.init = 16'hc088;
    LUT4 mux_1380_i22_3_lut (.A(n225[21]), .B(databus[21]), .C(n3446), 
         .Z(n3447[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i22_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i4 (.D(n5184[4]), .SP(n11908), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    CCU2D sub_126_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24411), .COUT(n24412), .S0(n225[13]), 
          .S1(n225[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_15.INIT0 = 16'h5555;
    defparam sub_126_add_2_15.INIT1 = 16'h5555;
    defparam sub_126_add_2_15.INJECT1_0 = "NO";
    defparam sub_126_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24410), .COUT(n24411), .S0(n225[11]), 
          .S1(n225[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_13.INIT0 = 16'h5555;
    defparam sub_126_add_2_13.INIT1 = 16'h5555;
    defparam sub_126_add_2_13.INJECT1_0 = "NO";
    defparam sub_126_add_2_13.INJECT1_1 = "NO";
    LUT4 mux_1380_i21_3_lut (.A(n225[20]), .B(databus[20]), .C(n3446), 
         .Z(n3447[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1380_i21_3_lut.init = 16'hcaca;
    CCU2D sub_126_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24409), .COUT(n24410), .S0(n225[9]), .S1(n225[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_11.INIT0 = 16'h5555;
    defparam sub_126_add_2_11.INIT1 = 16'h5555;
    defparam sub_126_add_2_11.INJECT1_0 = "NO";
    defparam sub_126_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_9 (.A0(\steps_reg[7] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24408), .COUT(n24409), .S0(n225[7]), .S1(n225[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_9.INIT0 = 16'h5555;
    defparam sub_126_add_2_9.INIT1 = 16'h5555;
    defparam sub_126_add_2_9.INJECT1_0 = "NO";
    defparam sub_126_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24407), .COUT(n24408), .S0(n225[5]), .S1(n225[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_7.INIT0 = 16'h5555;
    defparam sub_126_add_2_7.INIT1 = 16'h5555;
    defparam sub_126_add_2_7.INJECT1_0 = "NO";
    defparam sub_126_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24406), .COUT(n24407), .S0(n225[3]), .S1(n225[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_5.INIT0 = 16'h5555;
    defparam sub_126_add_2_5.INIT1 = 16'h5555;
    defparam sub_126_add_2_5.INJECT1_0 = "NO";
    defparam sub_126_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_126_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24405), .COUT(n24406), .S0(n225[1]), .S1(n225[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_3.INIT0 = 16'h5555;
    defparam sub_126_add_2_3.INIT1 = 16'h5555;
    defparam sub_126_add_2_3.INJECT1_0 = "NO";
    defparam sub_126_add_2_3.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_178 (.A(div_factor_reg[20]), .B(\register_addr[1] ), 
         .C(steps_reg[20]), .D(\register_addr[0] ), .Z(n26873)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_178.init = 16'hc088;
    CCU2D sub_126_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(step_clk), .C1(n21), .D1(prev_step_clk), 
          .COUT(n24405), .S1(n225[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_126_add_2_1.INIT0 = 16'h0000;
    defparam sub_126_add_2_1.INIT1 = 16'h5595;
    defparam sub_126_add_2_1.INJECT1_0 = "NO";
    defparam sub_126_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_179 (.A(div_factor_reg[21]), .B(\register_addr[1] ), 
         .C(steps_reg[21]), .D(\register_addr[0] ), .Z(n26877)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_179.init = 16'hc088;
    LUT4 i1_4_lut_adj_180 (.A(div_factor_reg[22]), .B(\register_addr[1] ), 
         .C(steps_reg[22]), .D(\register_addr[0] ), .Z(n26887)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_180.init = 16'hc088;
    LUT4 i1_4_lut_adj_181 (.A(div_factor_reg[23]), .B(\register_addr[1] ), 
         .C(steps_reg[23]), .D(\register_addr[0] ), .Z(n26886)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_181.init = 16'hc088;
    LUT4 i1_4_lut_adj_182 (.A(div_factor_reg[24]), .B(\register_addr[1] ), 
         .C(steps_reg[24]), .D(\register_addr[0] ), .Z(n26888)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_182.init = 16'hc088;
    LUT4 i1_4_lut_adj_183 (.A(div_factor_reg[25]), .B(\register_addr[1] ), 
         .C(steps_reg[25]), .D(\register_addr[0] ), .Z(n26889)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_183.init = 16'hc088;
    LUT4 i1_2_lut_4_lut (.A(n28917), .B(n29052), .C(n28898), .D(n30647), 
         .Z(n12444)) /* synthesis lut_function=(A (D)+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hff40;
    LUT4 i1_4_lut_adj_184 (.A(div_factor_reg[26]), .B(\register_addr[1] ), 
         .C(steps_reg[26]), .D(\register_addr[0] ), .Z(n26890)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_184.init = 16'hc088;
    LUT4 i1_4_lut_adj_185 (.A(div_factor_reg[27]), .B(\register_addr[1] ), 
         .C(steps_reg[27]), .D(\register_addr[0] ), .Z(n26891)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_185.init = 16'hc088;
    LUT4 i3843_3_lut (.A(prev_limit_latched), .B(n30647), .C(limit_latched), 
         .Z(n9604)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i3843_3_lut.init = 16'hdcdc;
    LUT4 i1_4_lut_adj_186 (.A(div_factor_reg[28]), .B(\register_addr[1] ), 
         .C(steps_reg[28]), .D(\register_addr[0] ), .Z(n26892)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_186.init = 16'hc088;
    LUT4 i1_4_lut_adj_187 (.A(div_factor_reg[29]), .B(\register_addr[1] ), 
         .C(steps_reg[29]), .D(\register_addr[0] ), .Z(n26893)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_187.init = 16'hc088;
    ClockDivider_U8 step_clk_gen (.GND_net(GND_net), .prev_step_clk(prev_step_clk), 
            .n21(n21), .step_clk(step_clk), .n28908(n28908), .n30647(n30647), 
            .n12(n12), .debug_c_c(debug_c_c), .div_factor_reg({div_factor_reg}), 
            .n28991(n28991)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U8
//

module ClockDivider_U8 (GND_net, prev_step_clk, n21, step_clk, n28908, 
            n30647, n12, debug_c_c, div_factor_reg, n28991) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input prev_step_clk;
    input n21;
    output step_clk;
    output n28908;
    input n30647;
    output n12;
    input debug_c_c;
    input [31:0]div_factor_reg;
    input n28991;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n24530;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n24531, n24529, n24528, n24155;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n24156, n24154, n24153, n24527, n24526, n24525, n24524, 
        n24152;
    wire [31:0]n40;
    
    wire n6844, n24151, n24150, n24149, n24148, n24147, n24146, 
        n24145, n28892, n14058, n24144, n24143, n24142, n6809, 
        n24141, n24140, n24139, n24138, n24137, n24356, n24355, 
        n24354, n24136, n6878, n24135, n24353, n24352, n24134, 
        n24351, n24350, n24349, n24133, n24132, n24348, n24347, 
        n24346, n24131, n24345, n24130, n24129, n24344, n24343, 
        n24342, n24128, n24341, n24127, n24126, n24125, n24124, 
        n24123, n24122, n24121, n24168, n24167, n24166, n24165, 
        n24164, n24163, n24162, n24161, n24160, n24159, n24158, 
        n24539, n24157, n24538, n24537, n24536, n24535, n24534, 
        n24533, n24532;
    
    CCU2D count_2168_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24530), .COUT(n24531), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2168_add_4_15.INJECT1_0 = "NO";
    defparam count_2168_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24529), .COUT(n24530), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2168_add_4_13.INJECT1_0 = "NO";
    defparam count_2168_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24528), .COUT(n24529), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2168_add_4_11.INJECT1_0 = "NO";
    defparam count_2168_add_4_11.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24155), .COUT(n24156));
    defparam sub_1710_add_2_7.INIT0 = 16'h5999;
    defparam sub_1710_add_2_7.INIT1 = 16'h5999;
    defparam sub_1710_add_2_7.INJECT1_0 = "NO";
    defparam sub_1710_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24154), .COUT(n24155));
    defparam sub_1710_add_2_5.INIT0 = 16'h5999;
    defparam sub_1710_add_2_5.INIT1 = 16'h5999;
    defparam sub_1710_add_2_5.INJECT1_0 = "NO";
    defparam sub_1710_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24153), .COUT(n24154));
    defparam sub_1710_add_2_3.INIT0 = 16'h5999;
    defparam sub_1710_add_2_3.INIT1 = 16'h5999;
    defparam sub_1710_add_2_3.INJECT1_0 = "NO";
    defparam sub_1710_add_2_3.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24527), .COUT(n24528), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2168_add_4_9.INJECT1_0 = "NO";
    defparam count_2168_add_4_9.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n24153));
    defparam sub_1710_add_2_1.INIT0 = 16'h0000;
    defparam sub_1710_add_2_1.INIT1 = 16'h5999;
    defparam sub_1710_add_2_1.INJECT1_0 = "NO";
    defparam sub_1710_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24526), .COUT(n24527), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2168_add_4_7.INJECT1_0 = "NO";
    defparam count_2168_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24525), .COUT(n24526), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2168_add_4_5.INJECT1_0 = "NO";
    defparam count_2168_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24524), .COUT(n24525), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2168_add_4_3.INJECT1_0 = "NO";
    defparam count_2168_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24524), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_1.INIT0 = 16'hF000;
    defparam count_2168_add_4_1.INIT1 = 16'h0555;
    defparam count_2168_add_4_1.INJECT1_0 = "NO";
    defparam count_2168_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_1712_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24152), .S1(n6844));
    defparam sub_1712_add_2_33.INIT0 = 16'h5999;
    defparam sub_1712_add_2_33.INIT1 = 16'h0000;
    defparam sub_1712_add_2_33.INJECT1_0 = "NO";
    defparam sub_1712_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1712_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24151), .COUT(n24152));
    defparam sub_1712_add_2_31.INIT0 = 16'h5999;
    defparam sub_1712_add_2_31.INIT1 = 16'h5999;
    defparam sub_1712_add_2_31.INJECT1_0 = "NO";
    defparam sub_1712_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1712_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24150), .COUT(n24151));
    defparam sub_1712_add_2_29.INIT0 = 16'h5999;
    defparam sub_1712_add_2_29.INIT1 = 16'h5999;
    defparam sub_1712_add_2_29.INJECT1_0 = "NO";
    defparam sub_1712_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1712_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24149), .COUT(n24150));
    defparam sub_1712_add_2_27.INIT0 = 16'h5999;
    defparam sub_1712_add_2_27.INIT1 = 16'h5999;
    defparam sub_1712_add_2_27.INJECT1_0 = "NO";
    defparam sub_1712_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1712_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24148), .COUT(n24149));
    defparam sub_1712_add_2_25.INIT0 = 16'h5999;
    defparam sub_1712_add_2_25.INIT1 = 16'h5999;
    defparam sub_1712_add_2_25.INJECT1_0 = "NO";
    defparam sub_1712_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1712_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24147), .COUT(n24148));
    defparam sub_1712_add_2_23.INIT0 = 16'h5999;
    defparam sub_1712_add_2_23.INIT1 = 16'h5999;
    defparam sub_1712_add_2_23.INJECT1_0 = "NO";
    defparam sub_1712_add_2_23.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_250 (.A(prev_step_clk), .B(n21), .C(step_clk), .Z(n28908)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam i2_3_lut_rep_250.init = 16'h4040;
    LUT4 i1_4_lut_4_lut (.A(prev_step_clk), .B(n21), .C(step_clk), .D(n30647), 
         .Z(n12)) /* synthesis lut_function=(!(A (C+(D))+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam i1_4_lut_4_lut.init = 16'h004a;
    CCU2D sub_1712_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24146), .COUT(n24147));
    defparam sub_1712_add_2_21.INIT0 = 16'h5999;
    defparam sub_1712_add_2_21.INIT1 = 16'h5999;
    defparam sub_1712_add_2_21.INJECT1_0 = "NO";
    defparam sub_1712_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1712_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24145), .COUT(n24146));
    defparam sub_1712_add_2_19.INIT0 = 16'h5999;
    defparam sub_1712_add_2_19.INIT1 = 16'h5999;
    defparam sub_1712_add_2_19.INJECT1_0 = "NO";
    defparam sub_1712_add_2_19.INJECT1_1 = "NO";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n28892), .PD(n14058), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    CCU2D sub_1712_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24144), .COUT(n24145));
    defparam sub_1712_add_2_17.INIT0 = 16'h5999;
    defparam sub_1712_add_2_17.INIT1 = 16'h5999;
    defparam sub_1712_add_2_17.INJECT1_0 = "NO";
    defparam sub_1712_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1712_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24143), .COUT(n24144));
    defparam sub_1712_add_2_15.INIT0 = 16'h5999;
    defparam sub_1712_add_2_15.INIT1 = 16'h5999;
    defparam sub_1712_add_2_15.INJECT1_0 = "NO";
    defparam sub_1712_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1712_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24142), .COUT(n24143));
    defparam sub_1712_add_2_13.INIT0 = 16'h5999;
    defparam sub_1712_add_2_13.INIT1 = 16'h5999;
    defparam sub_1712_add_2_13.INJECT1_0 = "NO";
    defparam sub_1712_add_2_13.INJECT1_1 = "NO";
    FD1S3IX clk_o_22 (.D(n6809), .CK(debug_c_c), .CD(n28991), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_1712_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24141), .COUT(n24142));
    defparam sub_1712_add_2_11.INIT0 = 16'h5999;
    defparam sub_1712_add_2_11.INIT1 = 16'h5999;
    defparam sub_1712_add_2_11.INJECT1_0 = "NO";
    defparam sub_1712_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1712_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24140), .COUT(n24141));
    defparam sub_1712_add_2_9.INIT0 = 16'h5999;
    defparam sub_1712_add_2_9.INIT1 = 16'h5999;
    defparam sub_1712_add_2_9.INJECT1_0 = "NO";
    defparam sub_1712_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1712_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24139), .COUT(n24140));
    defparam sub_1712_add_2_7.INIT0 = 16'h5999;
    defparam sub_1712_add_2_7.INIT1 = 16'h5999;
    defparam sub_1712_add_2_7.INJECT1_0 = "NO";
    defparam sub_1712_add_2_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    CCU2D sub_1712_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24138), .COUT(n24139));
    defparam sub_1712_add_2_5.INIT0 = 16'h5999;
    defparam sub_1712_add_2_5.INIT1 = 16'h5999;
    defparam sub_1712_add_2_5.INJECT1_0 = "NO";
    defparam sub_1712_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1712_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n24137), .COUT(n24138));
    defparam sub_1712_add_2_3.INIT0 = 16'h5999;
    defparam sub_1712_add_2_3.INIT1 = 16'h5999;
    defparam sub_1712_add_2_3.INJECT1_0 = "NO";
    defparam sub_1712_add_2_3.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    CCU2D sub_1712_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n24137));
    defparam sub_1712_add_2_1.INIT0 = 16'h0000;
    defparam sub_1712_add_2_1.INIT1 = 16'h5999;
    defparam sub_1712_add_2_1.INJECT1_0 = "NO";
    defparam sub_1712_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24356), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24355), .COUT(n24356), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24354), .COUT(n24355), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1713_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24136), .S1(n6878));
    defparam sub_1713_add_2_33.INIT0 = 16'hf555;
    defparam sub_1713_add_2_33.INIT1 = 16'h0000;
    defparam sub_1713_add_2_33.INJECT1_0 = "NO";
    defparam sub_1713_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1713_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24135), .COUT(n24136));
    defparam sub_1713_add_2_31.INIT0 = 16'hf555;
    defparam sub_1713_add_2_31.INIT1 = 16'hf555;
    defparam sub_1713_add_2_31.INJECT1_0 = "NO";
    defparam sub_1713_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24353), .COUT(n24354), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24352), .COUT(n24353), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1713_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24134), .COUT(n24135));
    defparam sub_1713_add_2_29.INIT0 = 16'hf555;
    defparam sub_1713_add_2_29.INIT1 = 16'hf555;
    defparam sub_1713_add_2_29.INJECT1_0 = "NO";
    defparam sub_1713_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24351), .COUT(n24352), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24350), .COUT(n24351), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24349), .COUT(n24350), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1713_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24133), .COUT(n24134));
    defparam sub_1713_add_2_27.INIT0 = 16'hf555;
    defparam sub_1713_add_2_27.INIT1 = 16'hf555;
    defparam sub_1713_add_2_27.INJECT1_0 = "NO";
    defparam sub_1713_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1713_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24132), .COUT(n24133));
    defparam sub_1713_add_2_25.INIT0 = 16'hf555;
    defparam sub_1713_add_2_25.INIT1 = 16'hf555;
    defparam sub_1713_add_2_25.INJECT1_0 = "NO";
    defparam sub_1713_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24348), .COUT(n24349), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    FD1S3IX count_2168__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i0.GSR = "ENABLED";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24347), .COUT(n24348), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24346), .COUT(n24347), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1713_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24131), .COUT(n24132));
    defparam sub_1713_add_2_23.INIT0 = 16'hf555;
    defparam sub_1713_add_2_23.INIT1 = 16'hf555;
    defparam sub_1713_add_2_23.INJECT1_0 = "NO";
    defparam sub_1713_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24345), .COUT(n24346), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    CCU2D sub_1713_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24130), .COUT(n24131));
    defparam sub_1713_add_2_21.INIT0 = 16'hf555;
    defparam sub_1713_add_2_21.INIT1 = 16'hf555;
    defparam sub_1713_add_2_21.INJECT1_0 = "NO";
    defparam sub_1713_add_2_21.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    CCU2D sub_1713_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24129), .COUT(n24130));
    defparam sub_1713_add_2_19.INIT0 = 16'hf555;
    defparam sub_1713_add_2_19.INIT1 = 16'hf555;
    defparam sub_1713_add_2_19.INJECT1_0 = "NO";
    defparam sub_1713_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24344), .COUT(n24345), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24343), .COUT(n24344), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24342), .COUT(n24343), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1713_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24128), .COUT(n24129));
    defparam sub_1713_add_2_17.INIT0 = 16'hf555;
    defparam sub_1713_add_2_17.INIT1 = 16'hf555;
    defparam sub_1713_add_2_17.INJECT1_0 = "NO";
    defparam sub_1713_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24341), .COUT(n24342), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    LUT4 i950_2_lut_rep_234 (.A(n6844), .B(n30647), .Z(n28892)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i950_2_lut_rep_234.init = 16'heeee;
    LUT4 i8437_2_lut_3_lut (.A(n6844), .B(n30647), .C(n6878), .Z(n14058)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i8437_2_lut_3_lut.init = 16'he0e0;
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24341), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1713_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24127), .COUT(n24128));
    defparam sub_1713_add_2_15.INIT0 = 16'hf555;
    defparam sub_1713_add_2_15.INIT1 = 16'hf555;
    defparam sub_1713_add_2_15.INJECT1_0 = "NO";
    defparam sub_1713_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1713_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24126), .COUT(n24127));
    defparam sub_1713_add_2_13.INIT0 = 16'hf555;
    defparam sub_1713_add_2_13.INIT1 = 16'hf555;
    defparam sub_1713_add_2_13.INJECT1_0 = "NO";
    defparam sub_1713_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1713_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24125), .COUT(n24126));
    defparam sub_1713_add_2_11.INIT0 = 16'hf555;
    defparam sub_1713_add_2_11.INIT1 = 16'hf555;
    defparam sub_1713_add_2_11.INJECT1_0 = "NO";
    defparam sub_1713_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1713_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24124), .COUT(n24125));
    defparam sub_1713_add_2_9.INIT0 = 16'hf555;
    defparam sub_1713_add_2_9.INIT1 = 16'hf555;
    defparam sub_1713_add_2_9.INJECT1_0 = "NO";
    defparam sub_1713_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1713_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24123), .COUT(n24124));
    defparam sub_1713_add_2_7.INIT0 = 16'hf555;
    defparam sub_1713_add_2_7.INIT1 = 16'hf555;
    defparam sub_1713_add_2_7.INJECT1_0 = "NO";
    defparam sub_1713_add_2_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    CCU2D sub_1713_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24122), .COUT(n24123));
    defparam sub_1713_add_2_5.INIT0 = 16'hf555;
    defparam sub_1713_add_2_5.INIT1 = 16'hf555;
    defparam sub_1713_add_2_5.INJECT1_0 = "NO";
    defparam sub_1713_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1713_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24121), .COUT(n24122));
    defparam sub_1713_add_2_3.INIT0 = 16'hf555;
    defparam sub_1713_add_2_3.INIT1 = 16'hf555;
    defparam sub_1713_add_2_3.INJECT1_0 = "NO";
    defparam sub_1713_add_2_3.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    CCU2D sub_1713_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n24121));
    defparam sub_1713_add_2_1.INIT0 = 16'h0000;
    defparam sub_1713_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1713_add_2_1.INJECT1_0 = "NO";
    defparam sub_1713_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1S3IX count_2168__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i1.GSR = "ENABLED";
    FD1S3IX count_2168__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i2.GSR = "ENABLED";
    FD1S3IX count_2168__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i3.GSR = "ENABLED";
    FD1S3IX count_2168__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i4.GSR = "ENABLED";
    FD1S3IX count_2168__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i5.GSR = "ENABLED";
    FD1S3IX count_2168__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i6.GSR = "ENABLED";
    FD1S3IX count_2168__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i7.GSR = "ENABLED";
    FD1S3IX count_2168__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i8.GSR = "ENABLED";
    FD1S3IX count_2168__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i9.GSR = "ENABLED";
    FD1S3IX count_2168__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i10.GSR = "ENABLED";
    FD1S3IX count_2168__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i11.GSR = "ENABLED";
    FD1S3IX count_2168__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i12.GSR = "ENABLED";
    FD1S3IX count_2168__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i13.GSR = "ENABLED";
    FD1S3IX count_2168__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i14.GSR = "ENABLED";
    FD1S3IX count_2168__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i15.GSR = "ENABLED";
    FD1S3IX count_2168__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i16.GSR = "ENABLED";
    FD1S3IX count_2168__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i17.GSR = "ENABLED";
    FD1S3IX count_2168__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i18.GSR = "ENABLED";
    FD1S3IX count_2168__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i19.GSR = "ENABLED";
    FD1S3IX count_2168__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i20.GSR = "ENABLED";
    FD1S3IX count_2168__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i21.GSR = "ENABLED";
    FD1S3IX count_2168__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i22.GSR = "ENABLED";
    FD1S3IX count_2168__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i23.GSR = "ENABLED";
    FD1S3IX count_2168__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i24.GSR = "ENABLED";
    FD1S3IX count_2168__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i25.GSR = "ENABLED";
    FD1S3IX count_2168__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i26.GSR = "ENABLED";
    FD1S3IX count_2168__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i27.GSR = "ENABLED";
    FD1S3IX count_2168__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i28.GSR = "ENABLED";
    FD1S3IX count_2168__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i29.GSR = "ENABLED";
    FD1S3IX count_2168__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i30.GSR = "ENABLED";
    FD1S3IX count_2168__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n28892), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168__i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n28892), .CD(n14058), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    CCU2D sub_1710_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24168), .S1(n6809));
    defparam sub_1710_add_2_33.INIT0 = 16'h5555;
    defparam sub_1710_add_2_33.INIT1 = 16'h0000;
    defparam sub_1710_add_2_33.INJECT1_0 = "NO";
    defparam sub_1710_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24167), .COUT(n24168));
    defparam sub_1710_add_2_31.INIT0 = 16'h5999;
    defparam sub_1710_add_2_31.INIT1 = 16'h5999;
    defparam sub_1710_add_2_31.INJECT1_0 = "NO";
    defparam sub_1710_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24166), .COUT(n24167));
    defparam sub_1710_add_2_29.INIT0 = 16'h5999;
    defparam sub_1710_add_2_29.INIT1 = 16'h5999;
    defparam sub_1710_add_2_29.INJECT1_0 = "NO";
    defparam sub_1710_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24165), .COUT(n24166));
    defparam sub_1710_add_2_27.INIT0 = 16'h5999;
    defparam sub_1710_add_2_27.INIT1 = 16'h5999;
    defparam sub_1710_add_2_27.INJECT1_0 = "NO";
    defparam sub_1710_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24164), .COUT(n24165));
    defparam sub_1710_add_2_25.INIT0 = 16'h5999;
    defparam sub_1710_add_2_25.INIT1 = 16'h5999;
    defparam sub_1710_add_2_25.INJECT1_0 = "NO";
    defparam sub_1710_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24163), .COUT(n24164));
    defparam sub_1710_add_2_23.INIT0 = 16'h5999;
    defparam sub_1710_add_2_23.INIT1 = 16'h5999;
    defparam sub_1710_add_2_23.INJECT1_0 = "NO";
    defparam sub_1710_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24162), .COUT(n24163));
    defparam sub_1710_add_2_21.INIT0 = 16'h5999;
    defparam sub_1710_add_2_21.INIT1 = 16'h5999;
    defparam sub_1710_add_2_21.INJECT1_0 = "NO";
    defparam sub_1710_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24161), .COUT(n24162));
    defparam sub_1710_add_2_19.INIT0 = 16'h5999;
    defparam sub_1710_add_2_19.INIT1 = 16'h5999;
    defparam sub_1710_add_2_19.INJECT1_0 = "NO";
    defparam sub_1710_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24160), .COUT(n24161));
    defparam sub_1710_add_2_17.INIT0 = 16'h5999;
    defparam sub_1710_add_2_17.INIT1 = 16'h5999;
    defparam sub_1710_add_2_17.INJECT1_0 = "NO";
    defparam sub_1710_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24159), .COUT(n24160));
    defparam sub_1710_add_2_15.INIT0 = 16'h5999;
    defparam sub_1710_add_2_15.INIT1 = 16'h5999;
    defparam sub_1710_add_2_15.INJECT1_0 = "NO";
    defparam sub_1710_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24158), .COUT(n24159));
    defparam sub_1710_add_2_13.INIT0 = 16'h5999;
    defparam sub_1710_add_2_13.INIT1 = 16'h5999;
    defparam sub_1710_add_2_13.INJECT1_0 = "NO";
    defparam sub_1710_add_2_13.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24539), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_33.INIT1 = 16'h0000;
    defparam count_2168_add_4_33.INJECT1_0 = "NO";
    defparam count_2168_add_4_33.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24157), .COUT(n24158));
    defparam sub_1710_add_2_11.INIT0 = 16'h5999;
    defparam sub_1710_add_2_11.INIT1 = 16'h5999;
    defparam sub_1710_add_2_11.INJECT1_0 = "NO";
    defparam sub_1710_add_2_11.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24538), .COUT(n24539), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2168_add_4_31.INJECT1_0 = "NO";
    defparam count_2168_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24537), .COUT(n24538), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2168_add_4_29.INJECT1_0 = "NO";
    defparam count_2168_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24536), .COUT(n24537), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2168_add_4_27.INJECT1_0 = "NO";
    defparam count_2168_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24535), .COUT(n24536), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2168_add_4_25.INJECT1_0 = "NO";
    defparam count_2168_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_1710_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n24156), .COUT(n24157));
    defparam sub_1710_add_2_9.INIT0 = 16'h5999;
    defparam sub_1710_add_2_9.INIT1 = 16'h5999;
    defparam sub_1710_add_2_9.INJECT1_0 = "NO";
    defparam sub_1710_add_2_9.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24534), .COUT(n24535), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2168_add_4_23.INJECT1_0 = "NO";
    defparam count_2168_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24533), .COUT(n24534), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2168_add_4_21.INJECT1_0 = "NO";
    defparam count_2168_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24532), .COUT(n24533), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2168_add_4_19.INJECT1_0 = "NO";
    defparam count_2168_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2168_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24531), .COUT(n24532), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2168_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2168_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2168_add_4_17.INJECT1_0 = "NO";
    defparam count_2168_add_4_17.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module RCPeripheral
//

module RCPeripheral (databus_out, n2, rw, databus, \read_value[9] , 
            n1, n29028, \read_value[9]_adj_1 , read_value, n28904, 
            n53, n2_adj_3, \read_value[8]_adj_4 , n1_adj_5, \read_value[8]_adj_6 , 
            \register_addr[0] , n4, \read_value[7]_adj_7 , n28928, \select[7] , 
            \read_value[7]_adj_8 , \read_value[7]_adj_9 , n28905, n30644, 
            read_value_adj_142, n64, n4_adj_18, n176, \read_value[6]_adj_19 , 
            \read_value[6]_adj_20 , \read_value[6]_adj_21 , n2_adj_22, 
            \read_value[17]_adj_23 , n1_adj_24, \read_value[17]_adj_25 , 
            n2_adj_26, \read_value[16]_adj_27 , n1_adj_28, \read_value[16]_adj_29 , 
            n2_adj_30, \read_value[15]_adj_31 , n1_adj_32, \read_value[15]_adj_33 , 
            n2_adj_34, \read_value[14]_adj_35 , n1_adj_36, \read_value[14]_adj_37 , 
            n4_adj_38, \read_value[5]_adj_39 , \read_value[5]_adj_40 , 
            \read_value[5]_adj_41 , n2_adj_42, \read_value[13]_adj_43 , 
            n1_adj_44, \register_addr[2] , \read_value[13]_adj_45 , n2_adj_46, 
            \read_value[31]_adj_47 , n1_adj_48, \read_value[31]_adj_49 , 
            n2_adj_50, \read_value[30]_adj_51 , n1_adj_52, n2_adj_53, 
            \read_value[12]_adj_54 , n1_adj_55, \read_value[12]_adj_56 , 
            \read_value[30]_adj_57 , \register_addr[1] , n2_adj_58, \read_value[29]_adj_59 , 
            n1_adj_60, \read_value[29]_adj_61 , n2_adj_62, \read_value[11]_adj_63 , 
            n1_adj_64, \read_value[11]_adj_65 , n2_adj_66, \read_value[10]_adj_67 , 
            n1_adj_68, \read_value[10]_adj_69 , n28955, read_size, \select[1] , 
            n29018, \sendcount[1] , n11253, \read_size[2]_adj_70 , n28937, 
            \reg_size[2] , n28946, \read_size[2]_adj_71 , n4_adj_72, 
            \read_value[4]_adj_73 , \read_value[4]_adj_74 , \read_value[4]_adj_75 , 
            n2_adj_76, \read_value[28]_adj_77 , n1_adj_78, \read_value[28]_adj_79 , 
            n2_adj_80, \read_value[27]_adj_81 , n1_adj_82, \read_value[27]_adj_83 , 
            n2_adj_84, n4_adj_85, \read_value[26]_adj_86 , n1_adj_87, 
            \read_value[3]_adj_88 , \read_value[26]_adj_89 , n2_adj_90, 
            \read_value[3]_adj_91 , \read_value[3]_adj_92 , \read_value[25]_adj_93 , 
            n1_adj_94, \read_value[25]_adj_95 , n2_adj_96, \read_value[24]_adj_97 , 
            n1_adj_98, \read_value[24]_adj_99 , n4_adj_100, \read_value[2]_adj_101 , 
            n2_adj_102, \read_value[2]_adj_103 , \read_value[2]_adj_104 , 
            \read_value[23]_adj_105 , n1_adj_106, \read_value[23]_adj_107 , 
            n2_adj_108, n1_adj_109, \read_value[22]_adj_110 , n1_adj_111, 
            \read_value[1]_adj_112 , n6, \read_value[22]_adj_113 , n2_adj_114, 
            \read_value[1]_adj_115 , \read_value[21]_adj_116 , n1_adj_117, 
            \read_value[21]_adj_118 , n2_adj_119, \read_value[20]_adj_120 , 
            n1_adj_121, \read_value[20]_adj_122 , n4_adj_123, \read_value[0]_adj_124 , 
            \read_value[0]_adj_125 , \read_value[0]_adj_126 , \read_size[2]_adj_127 , 
            \read_size[2]_adj_128 , n28927, n28974, \read_size[0]_adj_129 , 
            n9, \read_size[0]_adj_130 , \read_size[0]_adj_131 , n10, 
            \read_size[0]_adj_132 , \select[2] , n8, n2_adj_133, \read_value[19]_adj_134 , 
            n1_adj_135, n2_adj_136, \read_value[19]_adj_137 , \read_value[18]_adj_138 , 
            n1_adj_139, \read_value[18]_adj_140 , debug_c_c, n28893, 
            rc_ch8_c, GND_net, n27548, n27590, n11996, n24991, n27575, 
            rc_ch7_c, n11997, n27556, n24998, n1030, n1018, n27509, 
            n4_adj_141, rc_ch4_c, n54, n26690, n28888, n14053, n27569, 
            rc_ch3_c, n27527, n12104, n24988, n27582, n27640, n12804, 
            rc_ch2_c, n24993, n27493, n27638, n12807, rc_ch1_c, 
            n24976) /* synthesis syn_module_defined=1 */ ;
    input [31:0]databus_out;
    input n2;
    input rw;
    output [31:0]databus;
    input \read_value[9] ;
    input n1;
    input n29028;
    input \read_value[9]_adj_1 ;
    input [31:0]read_value;
    input n28904;
    input n53;
    input n2_adj_3;
    input \read_value[8]_adj_4 ;
    input n1_adj_5;
    input \read_value[8]_adj_6 ;
    input \register_addr[0] ;
    input n4;
    input \read_value[7]_adj_7 ;
    input n28928;
    input \select[7] ;
    input \read_value[7]_adj_8 ;
    input \read_value[7]_adj_9 ;
    input n28905;
    input n30644;
    input [7:0]read_value_adj_142;
    input n64;
    input n4_adj_18;
    input n176;
    input \read_value[6]_adj_19 ;
    input \read_value[6]_adj_20 ;
    input \read_value[6]_adj_21 ;
    input n2_adj_22;
    input \read_value[17]_adj_23 ;
    input n1_adj_24;
    input \read_value[17]_adj_25 ;
    input n2_adj_26;
    input \read_value[16]_adj_27 ;
    input n1_adj_28;
    input \read_value[16]_adj_29 ;
    input n2_adj_30;
    input \read_value[15]_adj_31 ;
    input n1_adj_32;
    input \read_value[15]_adj_33 ;
    input n2_adj_34;
    input \read_value[14]_adj_35 ;
    input n1_adj_36;
    input \read_value[14]_adj_37 ;
    input n4_adj_38;
    input \read_value[5]_adj_39 ;
    input \read_value[5]_adj_40 ;
    input \read_value[5]_adj_41 ;
    input n2_adj_42;
    input \read_value[13]_adj_43 ;
    input n1_adj_44;
    input \register_addr[2] ;
    input \read_value[13]_adj_45 ;
    input n2_adj_46;
    input \read_value[31]_adj_47 ;
    input n1_adj_48;
    input \read_value[31]_adj_49 ;
    input n2_adj_50;
    input \read_value[30]_adj_51 ;
    input n1_adj_52;
    input n2_adj_53;
    input \read_value[12]_adj_54 ;
    input n1_adj_55;
    input \read_value[12]_adj_56 ;
    input \read_value[30]_adj_57 ;
    input \register_addr[1] ;
    input n2_adj_58;
    input \read_value[29]_adj_59 ;
    input n1_adj_60;
    input \read_value[29]_adj_61 ;
    input n2_adj_62;
    input \read_value[11]_adj_63 ;
    input n1_adj_64;
    input \read_value[11]_adj_65 ;
    input n2_adj_66;
    input \read_value[10]_adj_67 ;
    input n1_adj_68;
    input \read_value[10]_adj_69 ;
    input n28955;
    input [2:0]read_size;
    input \select[1] ;
    output n29018;
    input \sendcount[1] ;
    output n11253;
    input \read_size[2]_adj_70 ;
    input n28937;
    output \reg_size[2] ;
    input n28946;
    input \read_size[2]_adj_71 ;
    input n4_adj_72;
    input \read_value[4]_adj_73 ;
    input \read_value[4]_adj_74 ;
    input \read_value[4]_adj_75 ;
    input n2_adj_76;
    input \read_value[28]_adj_77 ;
    input n1_adj_78;
    input \read_value[28]_adj_79 ;
    input n2_adj_80;
    input \read_value[27]_adj_81 ;
    input n1_adj_82;
    input \read_value[27]_adj_83 ;
    input n2_adj_84;
    input n4_adj_85;
    input \read_value[26]_adj_86 ;
    input n1_adj_87;
    input \read_value[3]_adj_88 ;
    input \read_value[26]_adj_89 ;
    input n2_adj_90;
    input \read_value[3]_adj_91 ;
    input \read_value[3]_adj_92 ;
    input \read_value[25]_adj_93 ;
    input n1_adj_94;
    input \read_value[25]_adj_95 ;
    input n2_adj_96;
    input \read_value[24]_adj_97 ;
    input n1_adj_98;
    input \read_value[24]_adj_99 ;
    input n4_adj_100;
    input \read_value[2]_adj_101 ;
    input n2_adj_102;
    input \read_value[2]_adj_103 ;
    input \read_value[2]_adj_104 ;
    input \read_value[23]_adj_105 ;
    input n1_adj_106;
    input \read_value[23]_adj_107 ;
    input n2_adj_108;
    input n1_adj_109;
    input \read_value[22]_adj_110 ;
    input n1_adj_111;
    input \read_value[1]_adj_112 ;
    input n6;
    input \read_value[22]_adj_113 ;
    input n2_adj_114;
    input \read_value[1]_adj_115 ;
    input \read_value[21]_adj_116 ;
    input n1_adj_117;
    input \read_value[21]_adj_118 ;
    input n2_adj_119;
    input \read_value[20]_adj_120 ;
    input n1_adj_121;
    input \read_value[20]_adj_122 ;
    input n4_adj_123;
    input \read_value[0]_adj_124 ;
    input \read_value[0]_adj_125 ;
    input \read_value[0]_adj_126 ;
    input \read_size[2]_adj_127 ;
    input \read_size[2]_adj_128 ;
    input n28927;
    input n28974;
    input \read_size[0]_adj_129 ;
    output n9;
    input \read_size[0]_adj_130 ;
    input \read_size[0]_adj_131 ;
    output n10;
    input \read_size[0]_adj_132 ;
    input \select[2] ;
    output n8;
    input n2_adj_133;
    input \read_value[19]_adj_134 ;
    input n1_adj_135;
    input n2_adj_136;
    input \read_value[19]_adj_137 ;
    input \read_value[18]_adj_138 ;
    input n1_adj_139;
    input \read_value[18]_adj_140 ;
    input debug_c_c;
    input n28893;
    input rc_ch8_c;
    input GND_net;
    output n27548;
    output n27590;
    input n11996;
    input n24991;
    output n27575;
    input rc_ch7_c;
    input n11997;
    output n27556;
    input n24998;
    output n1030;
    output n1018;
    output n27509;
    output n4_adj_141;
    input rc_ch4_c;
    output n54;
    input n26690;
    input n28888;
    input n14053;
    output n27569;
    input rc_ch3_c;
    output n27527;
    input n12104;
    input n24988;
    output n27582;
    output n27640;
    input n12804;
    input rc_ch2_c;
    input n24993;
    output n27493;
    output n27638;
    input n12807;
    input rc_ch1_c;
    input n24976;
    
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n10_c, n8_c, n10_adj_13, n8_adj_15;
    wire [7:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    wire [7:0]\register[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    
    wire n28627, n994;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    
    wire n28628;
    wire [7:0]\register[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    wire [7:0]\register[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    
    wire n28625;
    wire [7:0]\register[6] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    
    wire n28624, n13, n12, n6_c, n10_adj_19, n7, n28668, n28669, 
        n29029;
    wire [7:0]read_value_adj_246;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(212[12:22])
    
    wire n7_adj_20, n7_adj_21, n7_adj_23, n7_adj_24, n7_adj_25, n7_adj_26, 
        n28671, n28672, n13_adj_31, n12_adj_33, n6_adj_34;
    wire [2:0]read_size_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(213[12:21])
    
    wire n10_adj_36, n28791, n979, n28792, n28789, n28788, n10_adj_41, 
        n8_adj_43, n28800, n28799, n28017, n10_adj_47, n8_adj_49, 
        n28802, n1054, n28803, n10_adj_53, n8_adj_55, n1039, n28386, 
        n10_adj_59, n8_adj_61, n13_adj_65, n12_adj_67, n6_adj_68, 
        n10_adj_70, n10_adj_75, n8_adj_77, n28151, n28148, n28152, 
        n28385, n28147, n28146, n10_adj_81, n8_adj_83, n10_adj_87, 
        n8_adj_89, n10_adj_91, n8_adj_93, n28150, n28149, n10_adj_99, 
        n8_adj_101, n28383, n28382, n28037, n28038, n28019, n28040, 
        n28020, n28021, n28018, n28022, n1024, n28041, n10_adj_105, 
        n8_adj_107, n10_adj_111, n8_adj_113, n28805, n1009, n28388, 
        n28674, n28043, n28630, n28804, n28801, n7_adj_117, n6_adj_118, 
        n28793, n28790, n28794, n13_adj_121, n12_adj_123, n6_adj_124, 
        n10_adj_126, n28673, n28670, n10_adj_131, n8_adj_133, n28016, 
        n28629, n28626, n10_adj_137, n8_adj_139, n10_adj_143, n13_adj_145, 
        n12_adj_147, n6_adj_148, n8_adj_149, n10_adj_152, n10_adj_155, 
        n8_adj_159, n10_adj_165, n8_adj_167, n13_adj_171, n12_adj_173, 
        n6_adj_174, n10_adj_176, n10_adj_177, n8_adj_183, n10_adj_187, 
        n14, n10_adj_190, n7_adj_191, n8_adj_192, n12_adj_195, n10_adj_201, 
        n8_adj_204, n10_adj_208, n8_adj_210, n13_adj_214, n12_adj_216, 
        n6_adj_217, n10_adj_219, n28042, n28039, n10_adj_233, n8_adj_235, 
        n10_adj_237, n8_adj_241, n28387, n28384;
    
    LUT4 i5_4_lut (.A(databus_out[9]), .B(n10_c), .C(n2), .D(rw), .Z(databus[9])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut.init = 16'hfcfe;
    LUT4 i4_4_lut (.A(\read_value[9] ), .B(n8_c), .C(n1), .D(n29028), 
         .Z(n10_c)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut.init = 16'hfefc;
    LUT4 i2_4_lut (.A(\read_value[9]_adj_1 ), .B(read_value[9]), .C(n28904), 
         .D(n53), .Z(n8_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut.init = 16'heca0;
    LUT4 i5_4_lut_adj_62 (.A(databus_out[8]), .B(n10_adj_13), .C(n2_adj_3), 
         .D(rw), .Z(databus[8])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_62.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_63 (.A(\read_value[8]_adj_4 ), .B(n8_adj_15), .C(n1_adj_5), 
         .D(n29028), .Z(n10_adj_13)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_63.init = 16'hfefc;
    LUT4 i2_4_lut_adj_64 (.A(\read_value[8]_adj_6 ), .B(read_value[8]), 
         .C(n28904), .D(n53), .Z(n8_adj_15)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_64.init = 16'heca0;
    LUT4 n994_bdd_3_lut_21712 (.A(\register[2] [1]), .B(\register[3] [1]), 
         .C(\register_addr[0] ), .Z(n28627)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n994_bdd_3_lut_21712.init = 16'hcaca;
    LUT4 n994_bdd_3_lut_22313 (.A(n994), .B(\register_addr[0] ), .C(\register[1] [1]), 
         .Z(n28628)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n994_bdd_3_lut_22313.init = 16'he2e2;
    LUT4 register_addr_1__bdd_3_lut_21721 (.A(\register_addr[0] ), .B(\register[4] [1]), 
         .C(\register[5] [1]), .Z(n28625)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_21721.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_21720 (.A(\register[6] [1]), .B(\register_addr[0] ), 
         .Z(n28624)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_21720.init = 16'h2222;
    LUT4 i7_4_lut (.A(n13), .B(n4), .C(n12), .D(n6_c), .Z(databus[7])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i5_4_lut_adj_65 (.A(\read_value[7]_adj_7 ), .B(n10_adj_19), .C(n7), 
         .D(n28928), .Z(n13)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_65.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_21744 (.A(\register[6] [5]), .B(\register_addr[0] ), 
         .Z(n28668)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_21744.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut_21745 (.A(\register_addr[0] ), .B(\register[4] [5]), 
         .C(\register[5] [5]), .Z(n28669)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_21745.init = 16'he4e4;
    LUT4 i14_2_lut_rep_371 (.A(\select[7] ), .B(rw), .Z(n29029)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam i14_2_lut_rep_371.init = 16'h8888;
    LUT4 Select_3612_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_246[5]), 
         .Z(n7_adj_20)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3612_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3611_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_246[6]), 
         .Z(n7_adj_21)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3611_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3610_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_246[7]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3610_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3617_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_246[0]), 
         .Z(n7_adj_23)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3617_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3615_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_246[2]), 
         .Z(n7_adj_24)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3615_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3614_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_246[3]), 
         .Z(n7_adj_25)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3614_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3613_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_246[4]), 
         .Z(n7_adj_26)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3613_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 i4_4_lut_adj_66 (.A(\read_value[7]_adj_8 ), .B(\read_value[7]_adj_9 ), 
         .C(n28905), .D(n29028), .Z(n12)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_66.init = 16'heca0;
    LUT4 \register_1[[5__bdd_3_lut_22306  (.A(\register[2] [5]), .B(\register[3] [5]), 
         .C(\register_addr[0] ), .Z(n28671)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[5__bdd_3_lut_22306 .init = 16'hcaca;
    LUT4 \register_1[[5__bdd_2_lut_22307  (.A(\register[1] [5]), .B(\register_addr[0] ), 
         .Z(n28672)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[5__bdd_2_lut_22307 .init = 16'h8888;
    LUT4 Select_3610_i6_2_lut (.A(databus_out[7]), .B(n30644), .Z(n6_c)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3610_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_67 (.A(read_value[7]), .B(read_value_adj_142[7]), 
         .C(n53), .D(n64), .Z(n10_adj_19)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_67.init = 16'heca0;
    LUT4 i7_4_lut_adj_68 (.A(n13_adj_31), .B(n4_adj_18), .C(n12_adj_33), 
         .D(n6_adj_34), .Z(databus[6])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_68.init = 16'hfffe;
    FD1S3AX read_size_i1 (.D(n176), .CK(\select[7] ), .Q(read_size_c[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_size_i1.GSR = "ENABLED";
    LUT4 i5_4_lut_adj_69 (.A(\read_value[6]_adj_19 ), .B(n10_adj_36), .C(n7_adj_21), 
         .D(n28928), .Z(n13_adj_31)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_69.init = 16'hfefc;
    LUT4 i4_4_lut_adj_70 (.A(\read_value[6]_adj_20 ), .B(\read_value[6]_adj_21 ), 
         .C(n28905), .D(n29028), .Z(n12_adj_33)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_70.init = 16'heca0;
    LUT4 n979_bdd_3_lut_21783 (.A(\register[2] [0]), .B(\register[3] [0]), 
         .C(\register_addr[0] ), .Z(n28791)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n979_bdd_3_lut_21783.init = 16'hcaca;
    LUT4 Select_3611_i6_2_lut (.A(databus_out[6]), .B(rw), .Z(n6_adj_34)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3611_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_71 (.A(read_value[6]), .B(read_value_adj_142[6]), 
         .C(n53), .D(n64), .Z(n10_adj_36)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_71.init = 16'heca0;
    LUT4 n979_bdd_3_lut_22293 (.A(n979), .B(\register_addr[0] ), .C(\register[1] [0]), 
         .Z(n28792)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n979_bdd_3_lut_22293.init = 16'he2e2;
    LUT4 register_addr_1__bdd_3_lut_21790 (.A(\register_addr[0] ), .B(\register[4] [0]), 
         .C(\register[5] [0]), .Z(n28789)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_21790.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_21789 (.A(\register[6] [0]), .B(\register_addr[0] ), 
         .Z(n28788)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_21789.init = 16'h2222;
    LUT4 i5_4_lut_adj_72 (.A(databus_out[17]), .B(n10_adj_41), .C(n2_adj_22), 
         .D(rw), .Z(databus[17])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_72.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_73 (.A(\read_value[17]_adj_23 ), .B(n8_adj_43), .C(n1_adj_24), 
         .D(n29028), .Z(n10_adj_41)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_73.init = 16'hfefc;
    LUT4 i2_4_lut_adj_74 (.A(\read_value[17]_adj_25 ), .B(read_value[17]), 
         .C(n28904), .D(n53), .Z(n8_adj_43)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_74.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut (.A(\register_addr[0] ), .B(\register[4] [7]), 
         .C(\register[5] [7]), .Z(n28800)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut (.A(\register[6] [7]), .B(\register_addr[0] ), 
         .Z(n28799)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut_21484 (.A(\register_addr[0] ), .B(\register[4] [4]), 
         .C(\register[5] [4]), .Z(n28017)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_21484.init = 16'he4e4;
    LUT4 i5_4_lut_adj_75 (.A(databus_out[16]), .B(n10_adj_47), .C(n2_adj_26), 
         .D(rw), .Z(databus[16])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_75.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_76 (.A(\read_value[16]_adj_27 ), .B(n8_adj_49), .C(n1_adj_28), 
         .D(n29028), .Z(n10_adj_47)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_76.init = 16'hfefc;
    LUT4 n1054_bdd_3_lut_21793 (.A(\register[2] [7]), .B(\register[3] [7]), 
         .C(\register_addr[0] ), .Z(n28802)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1054_bdd_3_lut_21793.init = 16'hcaca;
    LUT4 i2_4_lut_adj_77 (.A(\read_value[16]_adj_29 ), .B(read_value[16]), 
         .C(n28904), .D(n53), .Z(n8_adj_49)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_77.init = 16'heca0;
    LUT4 n1054_bdd_3_lut_22283 (.A(n1054), .B(\register_addr[0] ), .C(\register[1] [7]), 
         .Z(n28803)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1054_bdd_3_lut_22283.init = 16'he2e2;
    LUT4 i5_4_lut_adj_78 (.A(databus_out[15]), .B(n10_adj_53), .C(n2_adj_30), 
         .D(rw), .Z(databus[15])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_78.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_79 (.A(\read_value[15]_adj_31 ), .B(n8_adj_55), .C(n1_adj_32), 
         .D(n29028), .Z(n10_adj_53)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_79.init = 16'hfefc;
    LUT4 n1039_bdd_3_lut_21756 (.A(n1039), .B(\register_addr[0] ), .C(\register[1] [6]), 
         .Z(n28386)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1039_bdd_3_lut_21756.init = 16'he2e2;
    LUT4 i2_4_lut_adj_80 (.A(\read_value[15]_adj_33 ), .B(read_value[15]), 
         .C(n28904), .D(n53), .Z(n8_adj_55)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_80.init = 16'heca0;
    LUT4 i5_4_lut_adj_81 (.A(databus_out[14]), .B(n10_adj_59), .C(n2_adj_34), 
         .D(rw), .Z(databus[14])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_81.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_82 (.A(\read_value[14]_adj_35 ), .B(n8_adj_61), .C(n1_adj_36), 
         .D(n29028), .Z(n10_adj_59)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_82.init = 16'hfefc;
    LUT4 i2_4_lut_adj_83 (.A(\read_value[14]_adj_37 ), .B(read_value[14]), 
         .C(n28904), .D(n53), .Z(n8_adj_61)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_83.init = 16'heca0;
    LUT4 i7_4_lut_adj_84 (.A(n13_adj_65), .B(n4_adj_38), .C(n12_adj_67), 
         .D(n6_adj_68), .Z(databus[5])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_84.init = 16'hfffe;
    LUT4 i5_4_lut_adj_85 (.A(\read_value[5]_adj_39 ), .B(n10_adj_70), .C(n7_adj_20), 
         .D(n28928), .Z(n13_adj_65)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_85.init = 16'hfefc;
    LUT4 i4_4_lut_adj_86 (.A(\read_value[5]_adj_40 ), .B(\read_value[5]_adj_41 ), 
         .C(n28905), .D(n29028), .Z(n12_adj_67)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_86.init = 16'heca0;
    LUT4 Select_3612_i6_2_lut (.A(databus_out[5]), .B(rw), .Z(n6_adj_68)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3612_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_87 (.A(read_value[5]), .B(read_value_adj_142[5]), 
         .C(n53), .D(n64), .Z(n10_adj_70)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_87.init = 16'heca0;
    LUT4 i5_4_lut_adj_88 (.A(databus_out[13]), .B(n10_adj_75), .C(n2_adj_42), 
         .D(rw), .Z(databus[13])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_88.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_89 (.A(\read_value[13]_adj_43 ), .B(n8_adj_77), .C(n1_adj_44), 
         .D(n29028), .Z(n10_adj_75)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_89.init = 16'hfefc;
    L6MUX21 i21541 (.D0(n28151), .D1(n28148), .SD(\register_addr[2] ), 
            .Z(n28152));
    LUT4 n1039_bdd_3_lut_21618 (.A(\register[2] [6]), .B(\register[3] [6]), 
         .C(\register_addr[0] ), .Z(n28385)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1039_bdd_3_lut_21618.init = 16'hcaca;
    LUT4 i2_4_lut_adj_90 (.A(\read_value[13]_adj_45 ), .B(read_value[13]), 
         .C(n28904), .D(n53), .Z(n8_adj_77)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_90.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_21615 (.A(\register_addr[0] ), .B(\register[4] [2]), 
         .C(\register[5] [2]), .Z(n28147)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_21615.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_21614 (.A(\register[6] [2]), .B(\register_addr[0] ), 
         .Z(n28146)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_21614.init = 16'h2222;
    LUT4 i5_4_lut_adj_91 (.A(databus_out[31]), .B(n10_adj_81), .C(n2_adj_46), 
         .D(rw), .Z(databus[31])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_91.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_92 (.A(\read_value[31]_adj_47 ), .B(n8_adj_83), .C(n1_adj_48), 
         .D(n29028), .Z(n10_adj_81)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_92.init = 16'hfefc;
    LUT4 i2_4_lut_adj_93 (.A(\read_value[31]_adj_49 ), .B(read_value[31]), 
         .C(n28904), .D(n53), .Z(n8_adj_83)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_93.init = 16'heca0;
    LUT4 i5_4_lut_adj_94 (.A(databus_out[30]), .B(n10_adj_87), .C(n2_adj_50), 
         .D(rw), .Z(databus[30])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_94.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_95 (.A(\read_value[30]_adj_51 ), .B(n8_adj_89), .C(n1_adj_52), 
         .D(n29028), .Z(n10_adj_87)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_95.init = 16'hfefc;
    LUT4 i5_4_lut_adj_96 (.A(databus_out[12]), .B(n10_adj_91), .C(n2_adj_53), 
         .D(rw), .Z(databus[12])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_96.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_97 (.A(\read_value[12]_adj_54 ), .B(n8_adj_93), .C(n1_adj_55), 
         .D(n29028), .Z(n10_adj_91)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_97.init = 16'hfefc;
    LUT4 i2_4_lut_adj_98 (.A(\read_value[12]_adj_56 ), .B(read_value[12]), 
         .C(n28904), .D(n53), .Z(n8_adj_93)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_98.init = 16'heca0;
    LUT4 i2_4_lut_adj_99 (.A(\read_value[30]_adj_57 ), .B(read_value[30]), 
         .C(n28904), .D(n53), .Z(n8_adj_89)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_99.init = 16'heca0;
    PFUMX i21539 (.BLUT(n28150), .ALUT(n28149), .C0(\register_addr[1] ), 
          .Z(n28151));
    LUT4 i5_4_lut_adj_100 (.A(databus_out[29]), .B(n10_adj_99), .C(n2_adj_58), 
         .D(rw), .Z(databus[29])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_100.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_101 (.A(\read_value[29]_adj_59 ), .B(n8_adj_101), 
         .C(n1_adj_60), .D(n29028), .Z(n10_adj_99)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_101.init = 16'hfefc;
    LUT4 i2_4_lut_adj_102 (.A(\read_value[29]_adj_61 ), .B(read_value[29]), 
         .C(n28904), .D(n53), .Z(n8_adj_101)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_102.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_21707 (.A(\register_addr[0] ), .B(\register[4] [6]), 
         .C(\register[5] [6]), .Z(n28383)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_21707.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_21706 (.A(\register[6] [6]), .B(\register_addr[0] ), 
         .Z(n28382)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_21706.init = 16'h2222;
    PFUMX i21536 (.BLUT(n28147), .ALUT(n28146), .C0(\register_addr[1] ), 
          .Z(n28148));
    LUT4 register_addr_1__bdd_2_lut_21520 (.A(\register[6] [3]), .B(\register_addr[0] ), 
         .Z(n28037)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_21520.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut_21521 (.A(\register_addr[0] ), .B(\register[4] [3]), 
         .C(\register[5] [3]), .Z(n28038)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_21521.init = 16'he4e4;
    LUT4 \register_1[[4__bdd_3_lut_21671  (.A(\register[2] [4]), .B(\register[3] [4]), 
         .C(\register_addr[0] ), .Z(n28019)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[4__bdd_3_lut_21671 .init = 16'hcaca;
    LUT4 n1024_bdd_3_lut_21497 (.A(\register[2] [3]), .B(\register[3] [3]), 
         .C(\register_addr[0] ), .Z(n28040)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1024_bdd_3_lut_21497.init = 16'hcaca;
    LUT4 \register_1[[4__bdd_2_lut_21672  (.A(\register[1] [4]), .B(\register_addr[0] ), 
         .Z(n28020)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[4__bdd_2_lut_21672 .init = 16'h8888;
    L6MUX21 i21481 (.D0(n28021), .D1(n28018), .SD(\register_addr[2] ), 
            .Z(n28022));
    LUT4 n1009_bdd_3_lut_21538 (.A(\register[2] [2]), .B(\register[3] [2]), 
         .C(\register_addr[0] ), .Z(n28149)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1009_bdd_3_lut_21538.init = 16'hcaca;
    LUT4 n1024_bdd_3_lut_21733 (.A(n1024), .B(\register_addr[0] ), .C(\register[1] [3]), 
         .Z(n28041)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1024_bdd_3_lut_21733.init = 16'he2e2;
    LUT4 i5_4_lut_adj_103 (.A(databus_out[11]), .B(n10_adj_105), .C(n2_adj_62), 
         .D(rw), .Z(databus[11])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_103.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_104 (.A(\read_value[11]_adj_63 ), .B(n8_adj_107), 
         .C(n1_adj_64), .D(n29028), .Z(n10_adj_105)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_104.init = 16'hfefc;
    LUT4 i2_4_lut_adj_105 (.A(\read_value[11]_adj_65 ), .B(read_value[11]), 
         .C(n28904), .D(n53), .Z(n8_adj_107)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_105.init = 16'heca0;
    LUT4 i5_4_lut_adj_106 (.A(databus_out[10]), .B(n10_adj_111), .C(n2_adj_66), 
         .D(rw), .Z(databus[10])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_106.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_107 (.A(\read_value[10]_adj_67 ), .B(n8_adj_113), 
         .C(n1_adj_68), .D(n29028), .Z(n10_adj_111)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_107.init = 16'hfefc;
    LUT4 i2_4_lut_adj_108 (.A(\read_value[10]_adj_69 ), .B(read_value[10]), 
         .C(n28904), .D(n53), .Z(n8_adj_113)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_108.init = 16'heca0;
    FD1S3IX read_value__i7 (.D(n28805), .CK(\select[7] ), .CD(n28955), 
            .Q(read_value_adj_246[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i7.GSR = "ENABLED";
    LUT4 n1009_bdd_3_lut_21566 (.A(n1009), .B(\register_addr[0] ), .C(\register[1] [2]), 
         .Z(n28150)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1009_bdd_3_lut_21566.init = 16'he2e2;
    LUT4 Select_3625_i1_2_lut_rep_360 (.A(read_size[1]), .B(\select[1] ), 
         .Z(n29018)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_3625_i1_2_lut_rep_360.init = 16'h8888;
    FD1S3IX read_value__i6 (.D(n28388), .CK(\select[7] ), .CD(n28955), 
            .Q(read_value_adj_246[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i6.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut (.A(read_size[1]), .B(\select[1] ), .C(\sendcount[1] ), 
         .Z(n11253)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7878;
    FD1S3IX read_value__i5 (.D(n28674), .CK(\select[7] ), .CD(n28955), 
            .Q(read_value_adj_246[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1S3IX read_value__i4 (.D(n28022), .CK(\select[7] ), .CD(n28955), 
            .Q(read_value_adj_246[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1S3IX read_value__i3 (.D(n28043), .CK(\select[7] ), .CD(n28955), 
            .Q(read_value_adj_246[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1S3IX read_value__i2 (.D(n28152), .CK(\select[7] ), .CD(n28955), 
            .Q(read_value_adj_246[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1S3IX read_value__i1 (.D(n28630), .CK(\select[7] ), .CD(n28955), 
            .Q(read_value_adj_246[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i1.GSR = "ENABLED";
    L6MUX21 i21796 (.D0(n28804), .D1(n28801), .SD(\register_addr[2] ), 
            .Z(n28805));
    PFUMX i21794 (.BLUT(n28803), .ALUT(n28802), .C0(\register_addr[1] ), 
          .Z(n28804));
    LUT4 i4_4_lut_adj_109 (.A(n7_adj_117), .B(\read_size[2]_adj_70 ), .C(n6_adj_118), 
         .D(n28937), .Z(\reg_size[2] )) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i4_4_lut_adj_109.init = 16'hfefa;
    PFUMX i21791 (.BLUT(n28800), .ALUT(n28799), .C0(\register_addr[1] ), 
          .Z(n28801));
    L6MUX21 i21786 (.D0(n28793), .D1(n28790), .SD(\register_addr[2] ), 
            .Z(n28794));
    PFUMX i21784 (.BLUT(n28792), .ALUT(n28791), .C0(\register_addr[1] ), 
          .Z(n28793));
    PFUMX i21781 (.BLUT(n28789), .ALUT(n28788), .C0(\register_addr[1] ), 
          .Z(n28790));
    LUT4 i2_4_lut_adj_110 (.A(n28946), .B(read_size[2]), .C(\read_size[2]_adj_71 ), 
         .D(\select[1] ), .Z(n7_adj_117)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_110.init = 16'heca0;
    LUT4 i7_4_lut_adj_111 (.A(n13_adj_121), .B(n4_adj_72), .C(n12_adj_123), 
         .D(n6_adj_124), .Z(databus[4])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_111.init = 16'hfffe;
    LUT4 i5_4_lut_adj_112 (.A(\read_value[4]_adj_73 ), .B(n10_adj_126), 
         .C(n7_adj_26), .D(n28928), .Z(n13_adj_121)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_112.init = 16'hfefc;
    LUT4 i4_4_lut_adj_113 (.A(\read_value[4]_adj_74 ), .B(\read_value[4]_adj_75 ), 
         .C(n28905), .D(n29028), .Z(n12_adj_123)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_113.init = 16'heca0;
    LUT4 Select_3613_i6_2_lut (.A(databus_out[4]), .B(n30644), .Z(n6_adj_124)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3613_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_114 (.A(read_value[4]), .B(read_value_adj_142[4]), 
         .C(n53), .D(n64), .Z(n10_adj_126)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_114.init = 16'heca0;
    L6MUX21 i21741 (.D0(n28673), .D1(n28670), .SD(\register_addr[2] ), 
            .Z(n28674));
    PFUMX i21739 (.BLUT(n28672), .ALUT(n28671), .C0(\register_addr[1] ), 
          .Z(n28673));
    LUT4 i5_4_lut_adj_115 (.A(databus_out[28]), .B(n10_adj_131), .C(n2_adj_76), 
         .D(rw), .Z(databus[28])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_115.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_116 (.A(\read_value[28]_adj_77 ), .B(n8_adj_133), 
         .C(n1_adj_78), .D(n29028), .Z(n10_adj_131)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_116.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_21483 (.A(\register[6] [4]), .B(\register_addr[0] ), 
         .Z(n28016)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_21483.init = 16'h2222;
    PFUMX i21737 (.BLUT(n28669), .ALUT(n28668), .C0(\register_addr[1] ), 
          .Z(n28670));
    L6MUX21 i21715 (.D0(n28629), .D1(n28626), .SD(\register_addr[2] ), 
            .Z(n28630));
    LUT4 i2_4_lut_adj_117 (.A(\read_value[28]_adj_79 ), .B(read_value[28]), 
         .C(n28904), .D(n53), .Z(n8_adj_133)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_117.init = 16'heca0;
    PFUMX i21713 (.BLUT(n28628), .ALUT(n28627), .C0(\register_addr[1] ), 
          .Z(n28629));
    PFUMX i21710 (.BLUT(n28625), .ALUT(n28624), .C0(\register_addr[1] ), 
          .Z(n28626));
    LUT4 i5_4_lut_adj_118 (.A(databus_out[27]), .B(n10_adj_137), .C(n2_adj_80), 
         .D(rw), .Z(databus[27])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_118.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_119 (.A(\read_value[27]_adj_81 ), .B(n8_adj_139), 
         .C(n1_adj_82), .D(n29028), .Z(n10_adj_137)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_119.init = 16'hfefc;
    LUT4 i2_4_lut_adj_120 (.A(\read_value[27]_adj_83 ), .B(read_value[27]), 
         .C(n28904), .D(n53), .Z(n8_adj_139)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_120.init = 16'heca0;
    LUT4 i5_4_lut_adj_121 (.A(databus_out[26]), .B(n10_adj_143), .C(n2_adj_84), 
         .D(rw), .Z(databus[26])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_121.init = 16'hfcfe;
    LUT4 i7_4_lut_adj_122 (.A(n13_adj_145), .B(n4_adj_85), .C(n12_adj_147), 
         .D(n6_adj_148), .Z(databus[3])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_122.init = 16'hfffe;
    LUT4 i4_4_lut_adj_123 (.A(\read_value[26]_adj_86 ), .B(n8_adj_149), 
         .C(n1_adj_87), .D(n29028), .Z(n10_adj_143)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_123.init = 16'hfefc;
    LUT4 i5_4_lut_adj_124 (.A(\read_value[3]_adj_88 ), .B(n10_adj_152), 
         .C(n7_adj_25), .D(n28928), .Z(n13_adj_145)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_124.init = 16'hfefc;
    LUT4 i2_4_lut_adj_125 (.A(\read_value[26]_adj_89 ), .B(read_value[26]), 
         .C(n28904), .D(n53), .Z(n8_adj_149)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_125.init = 16'heca0;
    LUT4 i5_4_lut_adj_126 (.A(databus_out[25]), .B(n10_adj_155), .C(n2_adj_90), 
         .D(rw), .Z(databus[25])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_126.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_127 (.A(\read_value[3]_adj_91 ), .B(\read_value[3]_adj_92 ), 
         .C(n28905), .D(n29028), .Z(n12_adj_147)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_127.init = 16'heca0;
    LUT4 i4_4_lut_adj_128 (.A(\read_value[25]_adj_93 ), .B(n8_adj_159), 
         .C(n1_adj_94), .D(n29028), .Z(n10_adj_155)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_128.init = 16'hfefc;
    LUT4 i2_4_lut_adj_129 (.A(\read_value[25]_adj_95 ), .B(read_value[25]), 
         .C(n28904), .D(n53), .Z(n8_adj_159)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_129.init = 16'heca0;
    LUT4 Select_3614_i6_2_lut (.A(databus_out[3]), .B(n30644), .Z(n6_adj_148)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3614_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_130 (.A(read_value[3]), .B(read_value_adj_142[3]), 
         .C(n53), .D(n64), .Z(n10_adj_152)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_130.init = 16'heca0;
    LUT4 i5_4_lut_adj_131 (.A(databus_out[24]), .B(n10_adj_165), .C(n2_adj_96), 
         .D(rw), .Z(databus[24])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_131.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_132 (.A(\read_value[24]_adj_97 ), .B(n8_adj_167), 
         .C(n1_adj_98), .D(n29028), .Z(n10_adj_165)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_132.init = 16'hfefc;
    LUT4 i2_4_lut_adj_133 (.A(\read_value[24]_adj_99 ), .B(read_value[24]), 
         .C(n28904), .D(n53), .Z(n8_adj_167)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_133.init = 16'heca0;
    LUT4 i7_4_lut_adj_134 (.A(n13_adj_171), .B(n4_adj_100), .C(n12_adj_173), 
         .D(n6_adj_174), .Z(databus[2])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_134.init = 16'hfffe;
    LUT4 i5_4_lut_adj_135 (.A(\read_value[2]_adj_101 ), .B(n10_adj_176), 
         .C(n7_adj_24), .D(n28928), .Z(n13_adj_171)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_135.init = 16'hfefc;
    LUT4 i5_4_lut_adj_136 (.A(databus_out[23]), .B(n10_adj_177), .C(n2_adj_102), 
         .D(rw), .Z(databus[23])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_136.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_137 (.A(\read_value[2]_adj_103 ), .B(\read_value[2]_adj_104 ), 
         .C(n28905), .D(n29028), .Z(n12_adj_173)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_137.init = 16'heca0;
    LUT4 Select_3615_i6_2_lut (.A(databus_out[2]), .B(n30644), .Z(n6_adj_174)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3615_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_138 (.A(read_value[2]), .B(read_value_adj_142[2]), 
         .C(n53), .D(n64), .Z(n10_adj_176)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_138.init = 16'heca0;
    LUT4 i4_4_lut_adj_139 (.A(\read_value[23]_adj_105 ), .B(n8_adj_183), 
         .C(n1_adj_106), .D(n29028), .Z(n10_adj_177)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_139.init = 16'hfefc;
    LUT4 i2_4_lut_adj_140 (.A(\read_value[23]_adj_107 ), .B(read_value[23]), 
         .C(n28904), .D(n53), .Z(n8_adj_183)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_140.init = 16'heca0;
    PFUMX i21479 (.BLUT(n28020), .ALUT(n28019), .C0(\register_addr[1] ), 
          .Z(n28021));
    LUT4 i5_4_lut_adj_141 (.A(databus_out[22]), .B(n10_adj_187), .C(n2_adj_108), 
         .D(rw), .Z(databus[22])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_141.init = 16'hfcfe;
    LUT4 i7_4_lut_adj_142 (.A(n1_adj_109), .B(n14), .C(n10_adj_190), .D(n7_adj_191), 
         .Z(databus[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_142.init = 16'hfffe;
    LUT4 i4_4_lut_adj_143 (.A(\read_value[22]_adj_110 ), .B(n8_adj_192), 
         .C(n1_adj_111), .D(n29028), .Z(n10_adj_187)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_143.init = 16'hfefc;
    LUT4 i6_4_lut (.A(\read_value[1]_adj_112 ), .B(n12_adj_195), .C(n6), 
         .D(n28904), .Z(n14)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut.init = 16'hfefc;
    LUT4 i2_4_lut_adj_144 (.A(\read_value[22]_adj_113 ), .B(read_value[22]), 
         .C(n28904), .D(n53), .Z(n8_adj_192)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_144.init = 16'heca0;
    LUT4 i2_4_lut_adj_145 (.A(read_value[1]), .B(read_value_adj_142[1]), 
         .C(n53), .D(n64), .Z(n10_adj_190)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_145.init = 16'heca0;
    LUT4 i5_4_lut_adj_146 (.A(databus_out[21]), .B(n10_adj_201), .C(n2_adj_114), 
         .D(rw), .Z(databus[21])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_146.init = 16'hfcfe;
    LUT4 Select_3616_i7_2_lut (.A(databus_out[1]), .B(n30644), .Z(n7_adj_191)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3616_i7_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_147 (.A(\read_value[1]_adj_115 ), .B(read_value_adj_246[1]), 
         .C(n28905), .D(n29029), .Z(n12_adj_195)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_147.init = 16'heca0;
    LUT4 i4_4_lut_adj_148 (.A(\read_value[21]_adj_116 ), .B(n8_adj_204), 
         .C(n1_adj_117), .D(n29028), .Z(n10_adj_201)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_148.init = 16'hfefc;
    LUT4 i2_4_lut_adj_149 (.A(\read_value[21]_adj_118 ), .B(read_value[21]), 
         .C(n28904), .D(n53), .Z(n8_adj_204)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_149.init = 16'heca0;
    LUT4 i5_4_lut_adj_150 (.A(databus_out[20]), .B(n10_adj_208), .C(n2_adj_119), 
         .D(rw), .Z(databus[20])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_150.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_151 (.A(\read_value[20]_adj_120 ), .B(n8_adj_210), 
         .C(n1_adj_121), .D(n29028), .Z(n10_adj_208)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_151.init = 16'hfefc;
    LUT4 i2_4_lut_adj_152 (.A(\read_value[20]_adj_122 ), .B(read_value[20]), 
         .C(n28904), .D(n53), .Z(n8_adj_210)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_152.init = 16'heca0;
    LUT4 i7_4_lut_adj_153 (.A(n13_adj_214), .B(n4_adj_123), .C(n12_adj_216), 
         .D(n6_adj_217), .Z(databus[0])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_153.init = 16'hfffe;
    LUT4 i5_4_lut_adj_154 (.A(\read_value[0]_adj_124 ), .B(n10_adj_219), 
         .C(n7_adj_23), .D(n28928), .Z(n13_adj_214)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_154.init = 16'hfefc;
    LUT4 i4_4_lut_adj_155 (.A(\read_value[0]_adj_125 ), .B(\read_value[0]_adj_126 ), 
         .C(n28905), .D(n29028), .Z(n12_adj_216)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_155.init = 16'heca0;
    LUT4 Select_3617_i6_2_lut (.A(databus_out[0]), .B(n30644), .Z(n6_adj_217)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3617_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_156 (.A(read_value[0]), .B(read_value_adj_142[0]), 
         .C(n53), .D(n64), .Z(n10_adj_219)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_156.init = 16'heca0;
    LUT4 i1_4_lut (.A(\read_size[2]_adj_127 ), .B(\read_size[2]_adj_128 ), 
         .C(n28927), .D(n28974), .Z(n6_adj_118)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut.init = 16'heca0;
    L6MUX21 i21500 (.D0(n28042), .D1(n28039), .SD(\register_addr[2] ), 
            .Z(n28043));
    PFUMX i21498 (.BLUT(n28041), .ALUT(n28040), .C0(\register_addr[1] ), 
          .Z(n28042));
    PFUMX i21495 (.BLUT(n28038), .ALUT(n28037), .C0(\register_addr[1] ), 
          .Z(n28039));
    PFUMX i21477 (.BLUT(n28017), .ALUT(n28016), .C0(\register_addr[1] ), 
          .Z(n28018));
    LUT4 i2_4_lut_adj_157 (.A(read_size[0]), .B(\read_size[0]_adj_129 ), 
         .C(\select[1] ), .D(n28937), .Z(n9)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_157.init = 16'heca0;
    LUT4 i3_4_lut (.A(n28946), .B(\read_size[0]_adj_130 ), .C(\read_size[0]_adj_131 ), 
         .D(n28974), .Z(n10)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut.init = 16'heca0;
    LUT4 i1_4_lut_adj_158 (.A(read_size_c[0]), .B(\read_size[0]_adj_132 ), 
         .C(\select[7] ), .D(\select[2] ), .Z(n8)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_158.init = 16'heca0;
    FD1S3IX read_value__i0 (.D(n28794), .CK(\select[7] ), .CD(n28955), 
            .Q(read_value_adj_246[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i5_4_lut_adj_159 (.A(databus_out[19]), .B(n10_adj_233), .C(n2_adj_133), 
         .D(rw), .Z(databus[19])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_159.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_160 (.A(\read_value[19]_adj_134 ), .B(n8_adj_235), 
         .C(n1_adj_135), .D(n29028), .Z(n10_adj_233)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_160.init = 16'hfefc;
    LUT4 i5_4_lut_adj_161 (.A(databus_out[18]), .B(n10_adj_237), .C(n2_adj_136), 
         .D(rw), .Z(databus[18])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_161.init = 16'hfcfe;
    LUT4 i2_4_lut_adj_162 (.A(\read_value[19]_adj_137 ), .B(read_value[19]), 
         .C(n28904), .D(n53), .Z(n8_adj_235)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_162.init = 16'heca0;
    LUT4 i4_4_lut_adj_163 (.A(\read_value[18]_adj_138 ), .B(n8_adj_241), 
         .C(n1_adj_139), .D(n29028), .Z(n10_adj_237)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_163.init = 16'hfefc;
    L6MUX21 i21621 (.D0(n28387), .D1(n28384), .SD(\register_addr[2] ), 
            .Z(n28388));
    PFUMX i21616 (.BLUT(n28383), .ALUT(n28382), .C0(\register_addr[1] ), 
          .Z(n28384));
    LUT4 i2_4_lut_adj_164 (.A(\read_value[18]_adj_140 ), .B(read_value[18]), 
         .C(n28904), .D(n53), .Z(n8_adj_241)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_164.init = 16'heca0;
    PFUMX i21619 (.BLUT(n28386), .ALUT(n28385), .C0(\register_addr[1] ), 
          .Z(n28387));
    PWMReceiver recv_ch8 (.debug_c_c(debug_c_c), .n28893(n28893), .rc_ch8_c(rc_ch8_c), 
            .GND_net(GND_net), .n27548(n27548), .n27590(n27590), .\register[6] ({\register[6] }), 
            .n11996(n11996), .n1054(n1054), .n24991(n24991)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(259[14] 263[36])
    PWMReceiver_U1 recv_ch7 (.GND_net(GND_net), .n27575(n27575), .debug_c_c(debug_c_c), 
            .n28893(n28893), .rc_ch7_c(rc_ch7_c), .\register[5] ({\register[5] }), 
            .n11997(n11997), .n27556(n27556), .n1039(n1039), .n24998(n24998)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(254[14] 258[36])
    PWMReceiver_U2 recv_ch4 (.n1030(n1030), .n1018(n1018), .n27509(n27509), 
            .n4(n4_adj_141), .debug_c_c(debug_c_c), .n28893(n28893), .rc_ch4_c(rc_ch4_c), 
            .GND_net(GND_net), .n54(n54), .n1024(n1024), .n26690(n26690), 
            .\register[4] ({\register[4] }), .n28888(n28888), .n14053(n14053)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(249[14] 253[36])
    PWMReceiver_U3 recv_ch3 (.n27569(n27569), .debug_c_c(debug_c_c), .n28893(n28893), 
            .rc_ch3_c(rc_ch3_c), .GND_net(GND_net), .n27527(n27527), .\register[3] ({\register[3] }), 
            .n12104(n12104), .n1009(n1009), .n24988(n24988)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(244[14] 248[36])
    PWMReceiver_U4 recv_ch2 (.GND_net(GND_net), .n27582(n27582), .n27640(n27640), 
            .n28893(n28893), .debug_c_c(debug_c_c), .\register[2] ({\register[2] }), 
            .n12804(n12804), .rc_ch2_c(rc_ch2_c), .n994(n994), .n24993(n24993)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(239[14] 243[36])
    PWMReceiver_U5 recv_ch1 (.n27493(n27493), .n27638(n27638), .debug_c_c(debug_c_c), 
            .n28893(n28893), .GND_net(GND_net), .\register[1] ({\register[1] }), 
            .n12807(n12807), .rc_ch1_c(rc_ch1_c), .n979(n979), .n24976(n24976)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(234[17] 238[36])
    
endmodule
//
// Verilog Description of module PWMReceiver
//

module PWMReceiver (debug_c_c, n28893, rc_ch8_c, GND_net, n27548, 
            n27590, \register[6] , n11996, n1054, n24991) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n28893;
    input rc_ch8_c;
    input GND_net;
    output n27548;
    output n27590;
    output [7:0]\register[6] ;
    input n11996;
    output n1054;
    input n24991;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    
    wire n4, n27011, n1048, n1060, n29053, n28943, n27078, n11729, 
        n28975, n28948, n27012, n28923, n28924, n20396, n23, n27289, 
        n126, n28947, n20505, n23984;
    wire [15:0]n116;
    
    wire n23983, n27077, n23982, n28902, n29022, n24872, n27001, 
        n14108;
    wire [7:0]n43;
    
    wire n26737;
    wire [7:0]n943;
    
    wire n5, n6, n25043, n11832, n27106, n128_adj_10, n23981, 
        n25046, n27108, n23980, n23979, n23978, n23977, n24272, 
        n24271, n24270, n24269;
    
    LUT4 i1_2_lut_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_49 (.A(count[6]), .B(count[7]), .C(count[5]), 
         .Z(n27011)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_3_lut_adj_49.init = 16'h8080;
    LUT4 i5_2_lut_rep_395 (.A(n1048), .B(n1060), .Z(n29053)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i5_2_lut_rep_395.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_50 (.A(n1048), .B(n1060), .C(n28943), .Z(n27078)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i1_2_lut_3_lut_adj_50.init = 16'hf4f4;
    LUT4 i1_2_lut_rep_317 (.A(count[9]), .B(n11729), .Z(n28975)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_317.init = 16'heeee;
    LUT4 i1_2_lut_rep_290_3_lut (.A(count[9]), .B(n11729), .C(count[8]), 
         .Z(n28948)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_290_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_265_3_lut_4_lut (.A(count[9]), .B(n11729), .C(n27012), 
         .D(count[8]), .Z(n28923)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_265_3_lut_4_lut.init = 16'hfffe;
    IFS1P3DX latched_in_45 (.D(rc_ch8_c), .SP(n28893), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1060));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1060), .SP(n28893), .CK(debug_c_c), .Q(n1048));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i20919_3_lut_4_lut (.A(n28924), .B(n20396), .C(n28975), .D(n23), 
         .Z(n27289)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[13:39])
    defparam i20919_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_289 (.A(n126), .B(count[1]), .C(count[0]), .Z(n28947)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i2_3_lut_rep_289.init = 16'h8080;
    LUT4 i1_2_lut_rep_266_4_lut (.A(n126), .B(count[1]), .C(count[0]), 
         .D(count[8]), .Z(n28924)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_266_4_lut.init = 16'h8000;
    LUT4 i14761_2_lut_4_lut (.A(n126), .B(count[1]), .C(count[0]), .D(n28948), 
         .Z(n20505)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i14761_2_lut_4_lut.init = 16'hff80;
    CCU2D add_1489_17 (.A0(count[15]), .B0(n29053), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n23984), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_17.INIT0 = 16'hd222;
    defparam add_1489_17.INIT1 = 16'h0000;
    defparam add_1489_17.INJECT1_0 = "NO";
    defparam add_1489_17.INJECT1_1 = "NO";
    CCU2D add_1489_15 (.A0(count[13]), .B0(n29053), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n29053), .C1(GND_net), .D1(GND_net), .CIN(n23983), 
          .COUT(n23984), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_15.INIT0 = 16'hd222;
    defparam add_1489_15.INIT1 = 16'hd222;
    defparam add_1489_15.INJECT1_0 = "NO";
    defparam add_1489_15.INJECT1_1 = "NO";
    LUT4 i21350_3_lut_3_lut_4_lut (.A(n27012), .B(n28948), .C(n20396), 
         .D(n28943), .Z(n27077)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i21350_3_lut_3_lut_4_lut.init = 16'h000e;
    CCU2D add_1489_13 (.A0(count[11]), .B0(n29053), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n29053), .C1(GND_net), .D1(GND_net), .CIN(n23982), 
          .COUT(n23983), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_13.INIT0 = 16'hd222;
    defparam add_1489_13.INIT1 = 16'hd222;
    defparam add_1489_13.INJECT1_0 = "NO";
    defparam add_1489_13.INJECT1_1 = "NO";
    LUT4 i21_3_lut_rep_244_4_lut (.A(count[8]), .B(n28947), .C(n28975), 
         .D(n20396), .Z(n28902)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i21_3_lut_rep_244_4_lut.init = 16'h00f8;
    LUT4 i1_2_lut_rep_364 (.A(n1060), .B(n1048), .Z(n29022)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_364.init = 16'hbbbb;
    LUT4 i21265_2_lut_3_lut (.A(n1060), .B(n1048), .C(n24872), .Z(n27548)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i21265_2_lut_3_lut.init = 16'h4040;
    LUT4 i21307_4_lut (.A(n27001), .B(n29053), .C(n28943), .D(n29022), 
         .Z(n27590)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i21307_4_lut.init = 16'h3031;
    LUT4 i3_4_lut (.A(n28948), .B(n27289), .C(n28947), .D(n27012), .Z(n27001)) /* synthesis lut_function=(!(A (B)+!A (B+!(C (D))))) */ ;
    defparam i3_4_lut.init = 16'h3222;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n11996), .PD(n14108), .CK(debug_c_c), 
            .Q(\register[6] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n11996), .PD(n14108), .CK(debug_c_c), 
            .Q(\register[6] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n11996), .PD(n14108), .CK(debug_c_c), 
            .Q(\register[6] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n11996), .PD(n14108), .CK(debug_c_c), 
            .Q(\register[6] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n11996), .PD(n14108), .CK(debug_c_c), 
            .Q(\register[6] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n11996), .PD(n14108), .CK(debug_c_c), 
            .Q(\register[6] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n11996), .PD(n14108), .CK(debug_c_c), 
            .Q(\register[6] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n11996), .PD(n14108), .CK(debug_c_c), 
            .Q(\register[6] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i3_4_lut_adj_51 (.A(n1048), .B(n28893), .C(n26737), .D(n20396), 
         .Z(n14108)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut_adj_51.init = 16'h0080;
    LUT4 i2_4_lut (.A(n28924), .B(n24872), .C(count[9]), .D(n1060), 
         .Z(n26737)) /* synthesis lut_function=(!(A ((D)+!B)+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i2_4_lut.init = 16'h00c8;
    LUT4 i14551_2_lut (.A(n943[1]), .B(n23), .Z(n43[1])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14551_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(count[8]), .B(n28975), .C(count[1]), .D(n126), 
         .Z(n23)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0222;
    LUT4 i14657_4_lut (.A(count[9]), .B(n11729), .C(n5), .D(n6), .Z(n20396)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;
    defparam i14657_4_lut.init = 16'heeec;
    LUT4 i1_4_lut_adj_52 (.A(count[7]), .B(count[4]), .C(count[5]), .D(n25043), 
         .Z(n5)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_4_lut_adj_52.init = 16'heaaa;
    LUT4 i2_2_lut (.A(count[8]), .B(count[6]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_53 (.A(count[1]), .B(count[3]), .C(count[2]), .D(count[0]), 
         .Z(n25043)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i3_4_lut_adj_53.init = 16'hfffe;
    LUT4 i3_4_lut_adj_54 (.A(count[12]), .B(n11832), .C(count[13]), .D(n27106), 
         .Z(n11729)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_54.init = 16'hfffe;
    LUT4 i1_2_lut (.A(count[15]), .B(count[14]), .Z(n11832)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_55 (.A(count[11]), .B(count[10]), .Z(n27106)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_55.init = 16'heeee;
    LUT4 i2_4_lut_adj_56 (.A(n28902), .B(n23), .C(n28923), .D(n20505), 
         .Z(n24872)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i2_4_lut_adj_56.init = 16'heefe;
    LUT4 i1_4_lut_adj_57 (.A(n128_adj_10), .B(n27011), .C(count[4]), .D(count[3]), 
         .Z(n27012)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_4_lut_adj_57.init = 16'hccc8;
    FD1P3IX valid_48 (.D(n27077), .SP(n24991), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1054));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_58 (.A(count[2]), .B(count[1]), .Z(n128_adj_10)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_58.init = 16'h8888;
    CCU2D add_1489_11 (.A0(count[9]), .B0(n29053), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n29053), .C1(GND_net), .D1(GND_net), .CIN(n23981), 
          .COUT(n23982), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_11.INIT0 = 16'hd222;
    defparam add_1489_11.INIT1 = 16'hd222;
    defparam add_1489_11.INJECT1_0 = "NO";
    defparam add_1489_11.INJECT1_1 = "NO";
    LUT4 i3_4_lut_adj_59 (.A(count[3]), .B(count[2]), .C(count[4]), .D(n27011), 
         .Z(n126)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i3_4_lut_adj_59.init = 16'h8000;
    LUT4 i14552_2_lut (.A(n943[2]), .B(n23), .Z(n43[2])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14552_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_60 (.A(n27106), .B(count[9]), .C(n25046), .D(n4), 
         .Z(n27108)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_60.init = 16'hfeee;
    LUT4 i14553_2_lut (.A(n943[3]), .B(n23), .Z(n43[3])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14553_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_61 (.A(count[3]), .B(count[4]), .C(n128_adj_10), 
         .D(count[5]), .Z(n25046)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_4_lut_adj_61.init = 16'hffec;
    CCU2D add_1489_9 (.A0(count[7]), .B0(n29053), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n29053), .C1(GND_net), .D1(GND_net), .CIN(n23980), 
          .COUT(n23981), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_9.INIT0 = 16'hd222;
    defparam add_1489_9.INIT1 = 16'hd222;
    defparam add_1489_9.INJECT1_0 = "NO";
    defparam add_1489_9.INJECT1_1 = "NO";
    CCU2D add_1489_7 (.A0(count[5]), .B0(n29053), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n29053), .C1(GND_net), .D1(GND_net), .CIN(n23979), 
          .COUT(n23980), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_7.INIT0 = 16'hd222;
    defparam add_1489_7.INIT1 = 16'hd222;
    defparam add_1489_7.INJECT1_0 = "NO";
    defparam add_1489_7.INJECT1_1 = "NO";
    LUT4 i14554_2_lut (.A(n943[4]), .B(n23), .Z(n43[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14554_2_lut.init = 16'h8888;
    CCU2D add_1489_5 (.A0(count[3]), .B0(n29053), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n29053), .C1(GND_net), .D1(GND_net), .CIN(n23978), 
          .COUT(n23979), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_5.INIT0 = 16'hd222;
    defparam add_1489_5.INIT1 = 16'hd222;
    defparam add_1489_5.INJECT1_0 = "NO";
    defparam add_1489_5.INJECT1_1 = "NO";
    LUT4 i14555_2_lut (.A(n943[5]), .B(n23), .Z(n43[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14555_2_lut.init = 16'h8888;
    LUT4 i14556_2_lut (.A(n943[6]), .B(n23), .Z(n43[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14556_2_lut.init = 16'h8888;
    LUT4 i14557_2_lut (.A(n943[7]), .B(n23), .Z(n43[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14557_2_lut.init = 16'h8888;
    CCU2D add_1489_3 (.A0(count[1]), .B0(n29053), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n29053), .C1(GND_net), .D1(GND_net), .CIN(n23977), 
          .COUT(n23978), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_3.INIT0 = 16'hd222;
    defparam add_1489_3.INIT1 = 16'hd222;
    defparam add_1489_3.INJECT1_0 = "NO";
    defparam add_1489_3.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24272), 
          .S0(n943[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_61_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_9.INIT1 = 16'h0000;
    defparam sub_61_add_2_9.INJECT1_0 = "NO";
    defparam sub_61_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24271), 
          .COUT(n24272), .S0(n943[5]), .S1(n943[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_61_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_61_add_2_7.INJECT1_0 = "NO";
    defparam sub_61_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24270), 
          .COUT(n24271), .S0(n943[3]), .S1(n943[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_61_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_61_add_2_5.INJECT1_0 = "NO";
    defparam sub_61_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24269), 
          .COUT(n24270), .S0(n943[1]), .S1(n943[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_61_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_61_add_2_3.INJECT1_0 = "NO";
    defparam sub_61_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24269), 
          .S1(n943[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_61_add_2_1.INIT0 = 16'hF000;
    defparam sub_61_add_2_1.INIT1 = 16'h5555;
    defparam sub_61_add_2_1.INJECT1_0 = "NO";
    defparam sub_61_add_2_1.INJECT1_1 = "NO";
    CCU2D add_1489_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n27078), .B1(n1060), .C1(count[0]), .D1(n1048), .COUT(n23977), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_1.INIT0 = 16'hF000;
    defparam add_1489_1.INIT1 = 16'ha565;
    defparam add_1489_1.INJECT1_0 = "NO";
    defparam add_1489_1.INJECT1_1 = "NO";
    LUT4 i14365_2_lut (.A(n943[0]), .B(n23), .Z(n43[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14365_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_rep_285 (.A(n11832), .B(count[13]), .C(count[12]), .D(n27108), 
         .Z(n28943)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_rep_285.init = 16'heaaa;
    
endmodule
//
// Verilog Description of module PWMReceiver_U1
//

module PWMReceiver_U1 (GND_net, n27575, debug_c_c, n28893, rc_ch7_c, 
            \register[5] , n11997, n27556, n1039, n24998) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n27575;
    input debug_c_c;
    input n28893;
    input rc_ch7_c;
    output [7:0]\register[5] ;
    input n11997;
    output n27556;
    output n1039;
    input n24998;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    
    wire n28950, n24723, n26958, n27254, n29024, n107, n28979, 
        n29000, n1033, n1045, n29031, n25135, n29059, n27110, 
        n23988;
    wire [15:0]n116;
    
    wire n23989, n23987, n24997, n27067, n29057, n27309, n54, 
        n28999, n23, n28976, n29058, n29012, n28938, n27343, n4, 
        n28926, n27071, n23986, n23985, n4_adj_6, n24876, n27111, 
        n28977, n10, n14087;
    wire [7:0]n43;
    
    wire n26735, n24;
    wire [7:0]n934;
    
    wire n27281, n4_adj_7, n4_adj_8, n24276, n24275, n24274, n24273, 
        n23992, n23991, n23990;
    
    LUT4 i20887_3_lut_4_lut (.A(count[8]), .B(n28950), .C(n24723), .D(n26958), 
         .Z(n27254)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i20887_3_lut_4_lut.init = 16'hfeee;
    LUT4 i1_2_lut_rep_366 (.A(count[4]), .B(count[5]), .Z(n29024)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_rep_366.init = 16'h8888;
    LUT4 i1_2_lut_rep_321_3_lut_4_lut (.A(count[4]), .B(count[5]), .C(n107), 
         .D(count[3]), .Z(n28979)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_rep_321_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_342_3_lut (.A(count[4]), .B(count[5]), .C(count[3]), 
         .Z(n29000)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_rep_342_3_lut.init = 16'h8080;
    LUT4 i5_2_lut_rep_373 (.A(n1033), .B(n1045), .Z(n29031)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i5_2_lut_rep_373.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n1033), .B(n1045), .C(n25135), .D(n29059), 
         .Z(n27110)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff4;
    CCU2D add_1485_9 (.A0(count[7]), .B0(n29031), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n29031), .C1(GND_net), .D1(GND_net), .CIN(n23988), 
          .COUT(n23989), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_9.INIT0 = 16'hd222;
    defparam add_1485_9.INIT1 = 16'hd222;
    defparam add_1485_9.INJECT1_0 = "NO";
    defparam add_1485_9.INJECT1_1 = "NO";
    CCU2D add_1485_7 (.A0(count[5]), .B0(n29031), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n29031), .C1(GND_net), .D1(GND_net), .CIN(n23987), 
          .COUT(n23988), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_7.INIT0 = 16'hd222;
    defparam add_1485_7.INIT1 = 16'hd222;
    defparam add_1485_7.INJECT1_0 = "NO";
    defparam add_1485_7.INJECT1_1 = "NO";
    LUT4 i21292_4_lut (.A(n29059), .B(n29031), .C(n25135), .D(n24997), 
         .Z(n27575)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i21292_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n27254), .B(n27067), .C(n29057), .D(n27309), .Z(n24997)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccce;
    LUT4 i20939_4_lut (.A(n54), .B(n28999), .C(n23), .D(n28976), .Z(n27309)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20939_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_399 (.A(count[11]), .B(count[10]), .Z(n29057)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_399.init = 16'heeee;
    LUT4 i1_2_lut_rep_292_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(count[9]), 
         .D(n28999), .Z(n28950)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_292_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_400 (.A(count[6]), .B(count[7]), .Z(n29058)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_400.init = 16'h8888;
    LUT4 i1_2_lut_rep_354_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n29012)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_354_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_401 (.A(count[15]), .B(count[14]), .Z(n29059)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_401.init = 16'heeee;
    LUT4 i2_3_lut_rep_341_4_lut (.A(count[15]), .B(count[14]), .C(count[12]), 
         .D(count[13]), .Z(n28999)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_341_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_280_3_lut (.A(count[15]), .B(count[14]), .C(n25135), 
         .Z(n28938)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_280_3_lut.init = 16'hfefe;
    LUT4 i20975_2_lut_rep_318 (.A(count[9]), .B(n27343), .Z(n28976)) /* synthesis lut_function=(A (B)) */ ;
    defparam i20975_2_lut_rep_318.init = 16'h8888;
    LUT4 i1_2_lut_4_lut (.A(n107), .B(count[0]), .C(n29012), .D(count[3]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_268_3_lut_4_lut (.A(n29057), .B(n28999), .C(count[8]), 
         .D(count[9]), .Z(n28926)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_268_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_35 (.A(n29057), .B(n28999), .C(n27343), 
         .D(count[9]), .Z(n27071)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_3_lut_4_lut_adj_35.init = 16'hfeee;
    LUT4 i2_3_lut_4_lut (.A(n107), .B(n29000), .C(n29058), .D(count[0]), 
         .Z(n26958)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_3_lut_4_lut.init = 16'h8000;
    IFS1P3DX latched_in_45 (.D(rc_ch7_c), .SP(n28893), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1045));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    CCU2D add_1485_5 (.A0(count[3]), .B0(n29031), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n29031), .C1(GND_net), .D1(GND_net), .CIN(n23986), 
          .COUT(n23987), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_5.INIT0 = 16'hd222;
    defparam add_1485_5.INIT1 = 16'hd222;
    defparam add_1485_5.INJECT1_0 = "NO";
    defparam add_1485_5.INJECT1_1 = "NO";
    FD1P3AX prev_in_46 (.D(n1045), .SP(n28893), .CK(debug_c_c), .Q(n1033));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    CCU2D add_1485_3 (.A0(count[1]), .B0(n29031), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n29031), .C1(GND_net), .D1(GND_net), .CIN(n23985), 
          .COUT(n23986), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_3.INIT0 = 16'hd222;
    defparam add_1485_3.INIT1 = 16'hd222;
    defparam add_1485_3.INJECT1_0 = "NO";
    defparam add_1485_3.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n29057), .D(n4_adj_6), 
         .Z(n25135)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i2_4_lut_adj_36 (.A(count[3]), .B(count[5]), .C(n107), .D(count[4]), 
         .Z(n24876)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_4_lut_adj_36.init = 16'hffec;
    LUT4 i1_2_lut (.A(count[1]), .B(count[2]), .Z(n107)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut.init = 16'h8888;
    CCU2D add_1485_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n27110), .B1(n1045), .C1(count[0]), .D1(n1033), .COUT(n23985), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_1.INIT0 = 16'hF000;
    defparam add_1485_1.INIT1 = 16'ha565;
    defparam add_1485_1.INJECT1_0 = "NO";
    defparam add_1485_1.INJECT1_1 = "NO";
    LUT4 i21348_3_lut_4_lut_4_lut (.A(n28938), .B(n27071), .C(n28926), 
         .D(n24723), .Z(n27111)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i21348_3_lut_4_lut_4_lut.init = 16'h1110;
    LUT4 i1_3_lut_4_lut (.A(count[8]), .B(n29058), .C(count[9]), .D(n24876), 
         .Z(n4_adj_6)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i3_3_lut_rep_319_4_lut (.A(count[8]), .B(n29058), .C(count[0]), 
         .D(n107), .Z(n28977)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_3_lut_rep_319_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_4_lut (.A(count[8]), .B(n29058), .C(n28979), .D(n28950), 
         .Z(n23)) /* synthesis lut_function=(!((B (C+(D))+!B (D))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_4_lut_4_lut.init = 16'h002a;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n28950), .C(n26958), 
         .D(n24723), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n11997), .PD(n14087), .CK(debug_c_c), 
            .Q(\register[5] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i21273_4_lut (.A(n54), .B(n27067), .C(n23), .D(n10), .Z(n27556)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i21273_4_lut.init = 16'h3332;
    LUT4 i3_4_lut (.A(n29059), .B(n26735), .C(n29057), .D(n28893), .Z(n14087)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut.init = 16'h0400;
    LUT4 i4_4_lut (.A(count[12]), .B(n24), .C(count[13]), .D(n27067), 
         .Z(n26735)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i4_4_lut.init = 16'h0004;
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n11997), .PD(n14087), .CK(debug_c_c), 
            .Q(\register[5] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n11997), .PD(n14087), .CK(debug_c_c), 
            .Q(\register[5] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n11997), .PD(n14087), .CK(debug_c_c), 
            .Q(\register[5] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n11997), .PD(n14087), .CK(debug_c_c), 
            .Q(\register[5] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n11997), .PD(n14087), .CK(debug_c_c), 
            .Q(\register[5] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n11997), .PD(n14087), .CK(debug_c_c), 
            .Q(\register[5] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n11997), .PD(n14087), .CK(debug_c_c), 
            .Q(\register[5] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    LUT4 i31_4_lut (.A(n29024), .B(n27343), .C(count[9]), .D(n4), .Z(n24)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i31_4_lut.init = 16'h3a30;
    LUT4 i1_2_lut_adj_37 (.A(n23), .B(n934[0]), .Z(n43[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_37.init = 16'h8888;
    LUT4 i20973_4_lut (.A(n27281), .B(count[6]), .C(n29024), .D(n4_adj_7), 
         .Z(n27343)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;
    defparam i20973_4_lut.init = 16'hffec;
    LUT4 i20911_4_lut (.A(count[1]), .B(count[0]), .C(count[3]), .D(count[2]), 
         .Z(n27281)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20911_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_38 (.A(count[7]), .B(count[8]), .Z(n4_adj_7)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_adj_38.init = 16'heeee;
    LUT4 i2_4_lut_adj_39 (.A(n29058), .B(n107), .C(count[5]), .D(n4_adj_8), 
         .Z(n24723)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_39.init = 16'ha080;
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_40 (.A(count[4]), .B(count[3]), .Z(n4_adj_8)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_adj_40.init = 16'heeee;
    LUT4 i1_2_lut_adj_41 (.A(n1045), .B(n1033), .Z(n27067)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_41.init = 16'hbbbb;
    LUT4 i21_4_lut (.A(n29000), .B(n27071), .C(n28950), .D(n28977), 
         .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[13:39])
    defparam i21_4_lut.init = 16'h3230;
    FD1P3IX valid_48 (.D(n27111), .SP(n24998), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1039));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    CCU2D sub_60_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24276), 
          .S0(n934[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_60_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_9.INIT1 = 16'h0000;
    defparam sub_60_add_2_9.INJECT1_0 = "NO";
    defparam sub_60_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_60_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24275), 
          .COUT(n24276), .S0(n934[5]), .S1(n934[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_60_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_60_add_2_7.INJECT1_0 = "NO";
    defparam sub_60_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_60_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24274), 
          .COUT(n24275), .S0(n934[3]), .S1(n934[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_60_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_60_add_2_5.INJECT1_0 = "NO";
    defparam sub_60_add_2_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_42 (.A(n23), .B(n934[1]), .Z(n43[1])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_42.init = 16'h8888;
    CCU2D sub_60_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24273), 
          .COUT(n24274), .S0(n934[1]), .S1(n934[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_60_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_60_add_2_3.INJECT1_0 = "NO";
    defparam sub_60_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_60_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24273), 
          .S1(n934[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_60_add_2_1.INIT0 = 16'hF000;
    defparam sub_60_add_2_1.INIT1 = 16'h5555;
    defparam sub_60_add_2_1.INJECT1_0 = "NO";
    defparam sub_60_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_43 (.A(n23), .B(n934[2]), .Z(n43[2])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_43.init = 16'h8888;
    LUT4 i1_2_lut_adj_44 (.A(n23), .B(n934[3]), .Z(n43[3])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_44.init = 16'h8888;
    CCU2D add_1485_17 (.A0(count[15]), .B0(n29031), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n23992), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_17.INIT0 = 16'hd222;
    defparam add_1485_17.INIT1 = 16'h0000;
    defparam add_1485_17.INJECT1_0 = "NO";
    defparam add_1485_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_45 (.A(n23), .B(n934[4]), .Z(n43[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_45.init = 16'h8888;
    CCU2D add_1485_15 (.A0(count[13]), .B0(n29031), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n29031), .C1(GND_net), .D1(GND_net), .CIN(n23991), 
          .COUT(n23992), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_15.INIT0 = 16'hd222;
    defparam add_1485_15.INIT1 = 16'hd222;
    defparam add_1485_15.INJECT1_0 = "NO";
    defparam add_1485_15.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_46 (.A(n23), .B(n934[5]), .Z(n43[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_46.init = 16'h8888;
    LUT4 i1_2_lut_adj_47 (.A(n23), .B(n934[6]), .Z(n43[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_47.init = 16'h8888;
    LUT4 i1_2_lut_adj_48 (.A(n23), .B(n934[7]), .Z(n43[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_48.init = 16'h8888;
    CCU2D add_1485_13 (.A0(count[11]), .B0(n29031), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n29031), .C1(GND_net), .D1(GND_net), .CIN(n23990), 
          .COUT(n23991), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_13.INIT0 = 16'hd222;
    defparam add_1485_13.INIT1 = 16'hd222;
    defparam add_1485_13.INJECT1_0 = "NO";
    defparam add_1485_13.INJECT1_1 = "NO";
    CCU2D add_1485_11 (.A0(count[9]), .B0(n29031), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n29031), .C1(GND_net), .D1(GND_net), .CIN(n23989), 
          .COUT(n23990), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_11.INIT0 = 16'hd222;
    defparam add_1485_11.INIT1 = 16'hd222;
    defparam add_1485_11.INJECT1_0 = "NO";
    defparam add_1485_11.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U2
//

module PWMReceiver_U2 (n1030, n1018, n27509, n4, debug_c_c, n28893, 
            rc_ch4_c, GND_net, n54, n1024, n26690, \register[4] , 
            n28888, n14053) /* synthesis syn_module_defined=1 */ ;
    output n1030;
    output n1018;
    output n27509;
    output n4;
    input debug_c_c;
    input n28893;
    input rc_ch4_c;
    input GND_net;
    output n54;
    output n1024;
    input n26690;
    output [7:0]\register[4] ;
    input n28888;
    input n14053;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n29032, n26691, n21798;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    wire [15:0]n4048;
    
    wire n29034, n29002, n25019, n5, n29035, n26954, n24681, n28983, 
        n26579, n23, n20535, n24671, n27269, n27268, n11877, n6, 
        n11770, n25172, n16546, n25024, n142, n4_adj_5, n57, n28982, 
        n27323;
    wire [15:0]n116;
    wire [7:0]n43;
    wire [7:0]n925;
    
    wire n24000, n23999, n23998, n24280, n23997, n24279, n23996, 
        n24278, n23995, n24277, n23994, n23993;
    
    LUT4 i1_2_lut_rep_374 (.A(n1030), .B(n1018), .Z(n29032)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut_rep_374.init = 16'hdddd;
    LUT4 i21226_4_lut_4_lut (.A(n1030), .B(n1018), .C(n26691), .D(n21798), 
         .Z(n27509)) /* synthesis lut_function=(!(A ((D)+!B)+!A (C (D)))) */ ;
    defparam i21226_4_lut_4_lut.init = 16'h05dd;
    LUT4 i1_2_lut_3_lut (.A(n1030), .B(n1018), .C(count[0]), .Z(n4048[0])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i1_2_lut_rep_376 (.A(count[4]), .B(count[5]), .Z(n29034)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_376.init = 16'h8888;
    LUT4 i1_2_lut_rep_344_3_lut (.A(count[4]), .B(count[5]), .C(count[1]), 
         .Z(n29002)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_344_3_lut.init = 16'h8080;
    LUT4 i1_3_lut_4_lut (.A(count[4]), .B(count[5]), .C(n25019), .D(count[7]), 
         .Z(n5)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i1_2_lut_rep_377 (.A(count[6]), .B(count[7]), .Z(n29035)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_377.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_26 (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n26954)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_3_lut_adj_26.init = 16'h8080;
    LUT4 i1_4_lut_4_lut (.A(n24681), .B(n28983), .C(n26579), .D(n23), 
         .Z(n4)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (D)) */ ;
    defparam i1_4_lut_4_lut.init = 16'hff02;
    LUT4 i2_3_lut_4_lut (.A(n24681), .B(n28983), .C(n21798), .D(n20535), 
         .Z(n24671)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h00e0;
    FD1P3AX prev_in_46 (.D(n1030), .SP(n28893), .CK(debug_c_c), .Q(n1018));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch4_c), .SP(n28893), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1030));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n27269), .B(n1018), .C(n27268), .D(n20535), .Z(n26691)) /* synthesis lut_function=(!(A (B)+!A (B ((D)+!C)))) */ ;
    defparam i1_4_lut.init = 16'h3373;
    LUT4 i20899_2_lut (.A(n54), .B(n23), .Z(n27269)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20899_2_lut.init = 16'heeee;
    LUT4 i14790_4_lut (.A(n5), .B(n11877), .C(count[9]), .D(n6), .Z(n20535)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i14790_4_lut.init = 16'hfcec;
    LUT4 i2_2_lut (.A(count[8]), .B(count[6]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3_4_lut (.A(count[3]), .B(count[1]), .C(count[2]), .D(count[0]), 
         .Z(n25019)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i21285_4_lut (.A(count[12]), .B(n11770), .C(n25172), .D(count[13]), 
         .Z(n21798)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B))) */ ;
    defparam i21285_4_lut.init = 16'h1333;
    LUT4 i2_4_lut (.A(n16546), .B(n25024), .C(count[9]), .D(n26954), 
         .Z(n25172)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i2_4_lut.init = 16'hfefa;
    LUT4 i2_4_lut_adj_27 (.A(count[3]), .B(count[5]), .C(n142), .D(count[4]), 
         .Z(n25024)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_4_lut_adj_27.init = 16'hffec;
    LUT4 i2_4_lut_adj_28 (.A(n29035), .B(n142), .C(count[5]), .D(n4_adj_5), 
         .Z(n24681)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_4_lut_adj_28.init = 16'ha080;
    LUT4 i1_2_lut (.A(count[3]), .B(count[4]), .Z(n4_adj_5)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_29 (.A(n11770), .B(count[12]), .C(count[13]), .D(n16546), 
         .Z(n11877)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut_adj_29.init = 16'hfffe;
    LUT4 i1_2_lut_adj_30 (.A(count[14]), .B(count[15]), .Z(n11770)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_adj_30.init = 16'heeee;
    LUT4 i1_2_lut_adj_31 (.A(count[10]), .B(count[11]), .Z(n16546)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_adj_31.init = 16'heeee;
    LUT4 i1_2_lut_adj_32 (.A(count[1]), .B(count[2]), .Z(n142)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_32.init = 16'h8888;
    LUT4 i3_4_lut_adj_33 (.A(n57), .B(n29035), .C(count[0]), .D(n29002), 
         .Z(n26579)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut_adj_33.init = 16'h8000;
    LUT4 i1_2_lut_adj_34 (.A(count[2]), .B(count[3]), .Z(n57)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_adj_34.init = 16'h8888;
    LUT4 i21_4_lut (.A(count[8]), .B(n20535), .C(n28982), .D(n26579), 
         .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[13:39])
    defparam i21_4_lut.init = 16'h3230;
    LUT4 i1_2_lut_rep_324 (.A(count[9]), .B(n11877), .Z(n28982)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i1_2_lut_rep_324.init = 16'heeee;
    LUT4 i1_2_lut_rep_325 (.A(count[9]), .B(n11877), .C(count[8]), .Z(n28983)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i1_2_lut_rep_325.init = 16'hfefe;
    LUT4 i15_4_lut_4_lut (.A(count[9]), .B(n11877), .C(count[8]), .D(n27323), 
         .Z(n23)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i15_4_lut_4_lut.init = 16'h0010;
    LUT4 i20953_3_lut_4_lut (.A(count[1]), .B(n29034), .C(n26954), .D(n57), 
         .Z(n27323)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20953_3_lut_4_lut.init = 16'h8000;
    FD1P3IX valid_48 (.D(n24671), .SP(n26690), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1024));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n28888), .PD(n14053), .CK(debug_c_c), 
            .Q(\register[4] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i20898_3_lut_4_lut (.A(count[8]), .B(n28982), .C(n24681), .D(n26579), 
         .Z(n27268)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i20898_3_lut_4_lut.init = 16'hfeee;
    LUT4 i14354_2_lut (.A(n925[0]), .B(n23), .Z(n43[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14354_2_lut.init = 16'h8888;
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n28888), .PD(n14053), .CK(debug_c_c), 
            .Q(\register[4] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n28888), .PD(n14053), .CK(debug_c_c), 
            .Q(\register[4] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n28888), .PD(n14053), .CK(debug_c_c), 
            .Q(\register[4] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n28888), .PD(n14053), .CK(debug_c_c), 
            .Q(\register[4] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n28888), .PD(n14053), .CK(debug_c_c), 
            .Q(\register[4] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n28888), .PD(n14053), .CK(debug_c_c), 
            .Q(\register[4] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n28888), .PD(n14053), .CK(debug_c_c), 
            .Q(\register[4] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    CCU2D add_1481_17 (.A0(n29032), .B0(count[15]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24000), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_17.INIT0 = 16'h7888;
    defparam add_1481_17.INIT1 = 16'h0000;
    defparam add_1481_17.INJECT1_0 = "NO";
    defparam add_1481_17.INJECT1_1 = "NO";
    CCU2D add_1481_15 (.A0(n29032), .B0(count[13]), .C0(GND_net), .D0(GND_net), 
          .A1(n29032), .B1(count[14]), .C1(GND_net), .D1(GND_net), .CIN(n23999), 
          .COUT(n24000), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_15.INIT0 = 16'h7888;
    defparam add_1481_15.INIT1 = 16'h7888;
    defparam add_1481_15.INJECT1_0 = "NO";
    defparam add_1481_15.INJECT1_1 = "NO";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    CCU2D add_1481_13 (.A0(n29032), .B0(count[11]), .C0(GND_net), .D0(GND_net), 
          .A1(n29032), .B1(count[12]), .C1(GND_net), .D1(GND_net), .CIN(n23998), 
          .COUT(n23999), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_13.INIT0 = 16'h7888;
    defparam add_1481_13.INIT1 = 16'h7888;
    defparam add_1481_13.INJECT1_0 = "NO";
    defparam add_1481_13.INJECT1_1 = "NO";
    CCU2D sub_59_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24280), 
          .S0(n925[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_59_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_9.INIT1 = 16'h0000;
    defparam sub_59_add_2_9.INJECT1_0 = "NO";
    defparam sub_59_add_2_9.INJECT1_1 = "NO";
    CCU2D add_1481_11 (.A0(n29032), .B0(count[9]), .C0(GND_net), .D0(GND_net), 
          .A1(n29032), .B1(count[10]), .C1(GND_net), .D1(GND_net), .CIN(n23997), 
          .COUT(n23998), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_11.INIT0 = 16'h7888;
    defparam add_1481_11.INIT1 = 16'h7888;
    defparam add_1481_11.INJECT1_0 = "NO";
    defparam add_1481_11.INJECT1_1 = "NO";
    CCU2D sub_59_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24279), 
          .COUT(n24280), .S0(n925[5]), .S1(n925[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_59_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_59_add_2_7.INJECT1_0 = "NO";
    defparam sub_59_add_2_7.INJECT1_1 = "NO";
    CCU2D add_1481_9 (.A0(n29032), .B0(count[7]), .C0(GND_net), .D0(GND_net), 
          .A1(n29032), .B1(count[8]), .C1(GND_net), .D1(GND_net), .CIN(n23996), 
          .COUT(n23997), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_9.INIT0 = 16'h7888;
    defparam add_1481_9.INIT1 = 16'h7888;
    defparam add_1481_9.INJECT1_0 = "NO";
    defparam add_1481_9.INJECT1_1 = "NO";
    CCU2D sub_59_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24278), 
          .COUT(n24279), .S0(n925[3]), .S1(n925[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_59_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_59_add_2_5.INJECT1_0 = "NO";
    defparam sub_59_add_2_5.INJECT1_1 = "NO";
    CCU2D add_1481_7 (.A0(count[5]), .B0(n29032), .C0(GND_net), .D0(GND_net), 
          .A1(n29032), .B1(count[6]), .C1(GND_net), .D1(GND_net), .CIN(n23995), 
          .COUT(n23996), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_7.INIT0 = 16'h7888;
    defparam add_1481_7.INIT1 = 16'h7888;
    defparam add_1481_7.INJECT1_0 = "NO";
    defparam add_1481_7.INJECT1_1 = "NO";
    CCU2D sub_59_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24277), 
          .COUT(n24278), .S0(n925[1]), .S1(n925[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_59_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_59_add_2_3.INJECT1_0 = "NO";
    defparam sub_59_add_2_3.INJECT1_1 = "NO";
    CCU2D add_1481_5 (.A0(n29032), .B0(count[3]), .C0(GND_net), .D0(GND_net), 
          .A1(n29032), .B1(count[4]), .C1(GND_net), .D1(GND_net), .CIN(n23994), 
          .COUT(n23995), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_5.INIT0 = 16'h7888;
    defparam add_1481_5.INIT1 = 16'h7888;
    defparam add_1481_5.INJECT1_0 = "NO";
    defparam add_1481_5.INJECT1_1 = "NO";
    CCU2D sub_59_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24277), 
          .S1(n925[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_59_add_2_1.INIT0 = 16'hF000;
    defparam sub_59_add_2_1.INIT1 = 16'h5555;
    defparam sub_59_add_2_1.INJECT1_0 = "NO";
    defparam sub_59_add_2_1.INJECT1_1 = "NO";
    CCU2D add_1481_3 (.A0(count[1]), .B0(n29032), .C0(GND_net), .D0(GND_net), 
          .A1(n29032), .B1(count[2]), .C1(GND_net), .D1(GND_net), .CIN(n23993), 
          .COUT(n23994), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_3.INIT0 = 16'h7888;
    defparam add_1481_3.INIT1 = 16'h7888;
    defparam add_1481_3.INJECT1_0 = "NO";
    defparam add_1481_3.INJECT1_1 = "NO";
    CCU2D add_1481_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n4048[0]), .B1(n1030), .C1(n1018), .D1(n21798), .COUT(n23993), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_1.INIT0 = 16'hF000;
    defparam add_1481_1.INIT1 = 16'h59aa;
    defparam add_1481_1.INJECT1_0 = "NO";
    defparam add_1481_1.INJECT1_1 = "NO";
    LUT4 i14544_2_lut (.A(n925[1]), .B(n23), .Z(n43[1])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14544_2_lut.init = 16'h8888;
    LUT4 i14546_2_lut (.A(n925[3]), .B(n23), .Z(n43[3])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14546_2_lut.init = 16'h8888;
    LUT4 i14547_2_lut (.A(n925[4]), .B(n23), .Z(n43[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14547_2_lut.init = 16'h8888;
    LUT4 i14545_2_lut (.A(n925[2]), .B(n23), .Z(n43[2])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14545_2_lut.init = 16'h8888;
    LUT4 i14548_2_lut (.A(n925[5]), .B(n23), .Z(n43[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14548_2_lut.init = 16'h8888;
    LUT4 i14549_2_lut (.A(n925[6]), .B(n23), .Z(n43[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14549_2_lut.init = 16'h8888;
    LUT4 i14550_2_lut (.A(n925[7]), .B(n23), .Z(n43[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14550_2_lut.init = 16'h8888;
    
endmodule
//
// Verilog Description of module PWMReceiver_U3
//

module PWMReceiver_U3 (n27569, debug_c_c, n28893, rc_ch3_c, GND_net, 
            n27527, \register[3] , n12104, n1009, n24988) /* synthesis syn_module_defined=1 */ ;
    output n27569;
    input debug_c_c;
    input n28893;
    input rc_ch3_c;
    input GND_net;
    output n27527;
    output [7:0]\register[3] ;
    input n12104;
    output n1009;
    input n24988;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    
    wire n29037, n4, n29038, n29003, n28954, n29039, n29040, n29005, 
        n29041, n29006, n29042, n29004, n26716, n29054, n28945, 
        n27073, n28930, n27265, n26715, n1003, n1015, n54, n26682, 
        n28984, n27114, n28986, n24847, n10, n26729, n14417, n24, 
        n11879, n25152, n25000;
    wire [7:0]n916;
    wire [7:0]n43;
    
    wire n24871, n6, n27104, n24008;
    wire [15:0]n116;
    
    wire n24007, n24006, n24005, n24004, n24003, n28985, n25049, 
        n24002, n27113, n24001, n24284, n24283, n24282, n24281;
    
    LUT4 i1_2_lut_rep_379 (.A(count[2]), .B(count[1]), .Z(n29037)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_379.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[4]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_380 (.A(count[11]), .B(count[10]), .Z(n29038)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_380.init = 16'heeee;
    LUT4 i1_2_lut_rep_296_3_lut_4_lut (.A(count[11]), .B(count[10]), .C(count[9]), 
         .D(n29003), .Z(n28954)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_296_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_381 (.A(count[15]), .B(count[14]), .Z(n29039)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_381.init = 16'heeee;
    LUT4 i2_3_lut_rep_345_4_lut (.A(count[15]), .B(count[14]), .C(count[13]), 
         .D(count[12]), .Z(n29003)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_345_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_382 (.A(count[7]), .B(count[6]), .Z(n29040)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_382.init = 16'h8888;
    LUT4 i1_2_lut_rep_347_3_lut (.A(count[7]), .B(count[6]), .C(count[8]), 
         .Z(n29005)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_347_3_lut.init = 16'h8080;
    LUT4 i2_3_lut_rep_383 (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n29041)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_rep_383.init = 16'h8080;
    LUT4 i1_2_lut_rep_348_4_lut (.A(count[2]), .B(count[3]), .C(count[1]), 
         .D(count[0]), .Z(n29006)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_348_4_lut.init = 16'h8000;
    LUT4 i14138_2_lut_rep_384 (.A(count[4]), .B(count[5]), .Z(n29042)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14138_2_lut_rep_384.init = 16'h8888;
    LUT4 i2_3_lut_rep_346_4_lut (.A(count[4]), .B(count[5]), .C(count[7]), 
         .D(count[6]), .Z(n29004)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_rep_346_4_lut.init = 16'h8000;
    LUT4 i21286_4_lut (.A(n26716), .B(n29054), .C(n28945), .D(n27073), 
         .Z(n27569)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i21286_4_lut.init = 16'h3031;
    LUT4 i3_4_lut (.A(n28930), .B(n29038), .C(n27265), .D(n26715), .Z(n26716)) /* synthesis lut_function=(!(A (B+!(D))+!A (B+!(C (D))))) */ ;
    defparam i3_4_lut.init = 16'h3200;
    LUT4 i5_2_lut_rep_396 (.A(n1003), .B(n1015), .Z(n29054)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i5_2_lut_rep_396.init = 16'h4444;
    LUT4 i3_4_lut_adj_18 (.A(n54), .B(n29003), .C(n26682), .D(n28984), 
         .Z(n26715)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut_adj_18.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_adj_19 (.A(n1003), .B(n1015), .C(n28945), .Z(n27114)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i1_2_lut_3_lut_adj_19.init = 16'hf4f4;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n28954), .C(n28986), 
         .D(n24847), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    IFS1P3DX latched_in_45 (.D(rc_ch3_c), .SP(n28893), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1015));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1015), .SP(n28893), .CK(debug_c_c), .Q(n1003));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i21244_4_lut (.A(n54), .B(n27073), .C(n26682), .D(n10), .Z(n27527)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i21244_4_lut.init = 16'h3323;
    LUT4 i3_4_lut_adj_20 (.A(n29039), .B(n26729), .C(n29038), .D(n28893), 
         .Z(n14417)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut_adj_20.init = 16'h0400;
    LUT4 i4_4_lut (.A(count[13]), .B(n24), .C(count[12]), .D(n27073), 
         .Z(n26729)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i4_4_lut.init = 16'h0004;
    LUT4 i20815_4_lut_rep_287 (.A(n29039), .B(count[13]), .C(count[12]), 
         .D(n11879), .Z(n28945)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i20815_4_lut_rep_287.init = 16'heaaa;
    LUT4 i31_3_lut (.A(n25152), .B(n25000), .C(count[9]), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i31_3_lut.init = 16'h3a3a;
    LUT4 i14349_2_lut (.A(n916[0]), .B(n26682), .Z(n43[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14349_2_lut.init = 16'h2222;
    LUT4 i1_4_lut (.A(n28954), .B(count[8]), .C(n29041), .D(n29004), 
         .Z(n26682)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfbbb;
    LUT4 i3_4_lut_adj_21 (.A(n24871), .B(n6), .C(count[6]), .D(n29042), 
         .Z(n25000)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_21.init = 16'hfefc;
    LUT4 i3_4_lut_adj_22 (.A(count[0]), .B(count[3]), .C(count[2]), .D(count[1]), 
         .Z(n24871)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_22.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[8]), .B(count[7]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1_2_lut (.A(n1015), .B(n1003), .Z(n27073)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i2_4_lut (.A(n29040), .B(count[3]), .C(count[5]), .D(n4), .Z(n24847)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_4_lut.init = 16'ha080;
    LUT4 i14828_2_lut_rep_326 (.A(n25000), .B(count[9]), .Z(n28984)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14828_2_lut_rep_326.init = 16'h8888;
    LUT4 i1_2_lut_rep_272_3_lut_4_lut (.A(n29038), .B(n29003), .C(count[8]), 
         .D(count[9]), .Z(n28930)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_272_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n29038), .B(n29003), .C(count[9]), .D(n25000), 
         .Z(n27104)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfeee;
    CCU2D add_1477_17 (.A0(count[15]), .B0(n29054), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24008), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_17.INIT0 = 16'hd222;
    defparam add_1477_17.INIT1 = 16'h0000;
    defparam add_1477_17.INJECT1_0 = "NO";
    defparam add_1477_17.INJECT1_1 = "NO";
    CCU2D add_1477_15 (.A0(count[13]), .B0(n29054), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n29054), .C1(GND_net), .D1(GND_net), .CIN(n24007), 
          .COUT(n24008), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_15.INIT0 = 16'hd222;
    defparam add_1477_15.INIT1 = 16'hd222;
    defparam add_1477_15.INJECT1_0 = "NO";
    defparam add_1477_15.INJECT1_1 = "NO";
    CCU2D add_1477_13 (.A0(count[11]), .B0(n29054), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n29054), .C1(GND_net), .D1(GND_net), .CIN(n24006), 
          .COUT(n24007), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_13.INIT0 = 16'hd222;
    defparam add_1477_13.INIT1 = 16'hd222;
    defparam add_1477_13.INJECT1_0 = "NO";
    defparam add_1477_13.INJECT1_1 = "NO";
    CCU2D add_1477_11 (.A0(count[9]), .B0(n29054), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n29054), .C1(GND_net), .D1(GND_net), .CIN(n24005), 
          .COUT(n24006), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_11.INIT0 = 16'hd222;
    defparam add_1477_11.INIT1 = 16'hd222;
    defparam add_1477_11.INJECT1_0 = "NO";
    defparam add_1477_11.INJECT1_1 = "NO";
    CCU2D add_1477_9 (.A0(count[7]), .B0(n29054), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n29054), .C1(GND_net), .D1(GND_net), .CIN(n24004), 
          .COUT(n24005), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_9.INIT0 = 16'hd222;
    defparam add_1477_9.INIT1 = 16'hd222;
    defparam add_1477_9.INJECT1_0 = "NO";
    defparam add_1477_9.INJECT1_1 = "NO";
    CCU2D add_1477_7 (.A0(count[5]), .B0(n29054), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n29054), .C1(GND_net), .D1(GND_net), .CIN(n24003), 
          .COUT(n24004), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_7.INIT0 = 16'hd222;
    defparam add_1477_7.INIT1 = 16'hd222;
    defparam add_1477_7.INJECT1_0 = "NO";
    defparam add_1477_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_327_4_lut (.A(count[12]), .B(n29039), .C(count[13]), 
         .D(n29038), .Z(n28985)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_327_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_328_4_lut (.A(count[6]), .B(count[7]), .C(n29042), 
         .D(n29006), .Z(n28986)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_328_4_lut.init = 16'h8000;
    LUT4 i3_3_lut_4_lut (.A(count[8]), .B(n29040), .C(n29006), .D(n29042), 
         .Z(n25152)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_23 (.A(count[0]), .B(n29041), .C(n24847), 
         .D(n29004), .Z(n27265)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_23.init = 16'h8000;
    LUT4 n25152_bdd_4_lut_21686 (.A(n25152), .B(count[9]), .C(n25000), 
         .D(n28985), .Z(n54)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A ((C+(D))+!B))) */ ;
    defparam n25152_bdd_4_lut_21686.init = 16'h002e;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n12104), .PD(n14417), .CK(debug_c_c), 
            .Q(\register[3] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i14543_2_lut (.A(n916[7]), .B(n26682), .Z(n43[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14543_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_24 (.A(n29038), .B(n25049), .C(count[9]), .D(n29005), 
         .Z(n11879)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i2_4_lut_adj_24.init = 16'hfefa;
    LUT4 i2_4_lut_adj_25 (.A(count[3]), .B(count[5]), .C(n29037), .D(count[4]), 
         .Z(n25049)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_4_lut_adj_25.init = 16'hffec;
    CCU2D add_1477_5 (.A0(count[3]), .B0(n29054), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n29054), .C1(GND_net), .D1(GND_net), .CIN(n24002), 
          .COUT(n24003), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_5.INIT0 = 16'hd222;
    defparam add_1477_5.INIT1 = 16'hd222;
    defparam add_1477_5.INJECT1_0 = "NO";
    defparam add_1477_5.INJECT1_1 = "NO";
    LUT4 i14542_2_lut (.A(n916[6]), .B(n26682), .Z(n43[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14542_2_lut.init = 16'h2222;
    LUT4 i14541_2_lut (.A(n916[5]), .B(n26682), .Z(n43[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14541_2_lut.init = 16'h2222;
    LUT4 i14540_2_lut (.A(n916[4]), .B(n26682), .Z(n43[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14540_2_lut.init = 16'h2222;
    LUT4 i14539_2_lut (.A(n916[3]), .B(n26682), .Z(n43[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14539_2_lut.init = 16'h2222;
    LUT4 i14538_2_lut (.A(n916[2]), .B(n26682), .Z(n43[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14538_2_lut.init = 16'h2222;
    LUT4 i21289_3_lut_4_lut_4_lut (.A(n28945), .B(n27104), .C(n28930), 
         .D(n24847), .Z(n27113)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i21289_3_lut_4_lut_4_lut.init = 16'h1110;
    LUT4 i14537_2_lut (.A(n916[1]), .B(n26682), .Z(n43[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14537_2_lut.init = 16'h2222;
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    CCU2D add_1477_3 (.A0(count[1]), .B0(n29054), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n29054), .C1(GND_net), .D1(GND_net), .CIN(n24001), 
          .COUT(n24002), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_3.INIT0 = 16'hd222;
    defparam add_1477_3.INIT1 = 16'hd222;
    defparam add_1477_3.INJECT1_0 = "NO";
    defparam add_1477_3.INJECT1_1 = "NO";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n12104), .PD(n14417), .CK(debug_c_c), 
            .Q(\register[3] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    CCU2D add_1477_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n27114), .B1(n1015), .C1(count[0]), .D1(n1003), .COUT(n24001), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_1.INIT0 = 16'hF000;
    defparam add_1477_1.INIT1 = 16'ha565;
    defparam add_1477_1.INJECT1_0 = "NO";
    defparam add_1477_1.INJECT1_1 = "NO";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n12104), .PD(n14417), .CK(debug_c_c), 
            .Q(\register[3] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n12104), .PD(n14417), .CK(debug_c_c), 
            .Q(\register[3] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n12104), .PD(n14417), .CK(debug_c_c), 
            .Q(\register[3] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n12104), .PD(n14417), .CK(debug_c_c), 
            .Q(\register[3] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n12104), .PD(n14417), .CK(debug_c_c), 
            .Q(\register[3] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n12104), .PD(n14417), .CK(debug_c_c), 
            .Q(\register[3] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D sub_58_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24284), 
          .S0(n916[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_58_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_9.INIT1 = 16'h0000;
    defparam sub_58_add_2_9.INJECT1_0 = "NO";
    defparam sub_58_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24283), 
          .COUT(n24284), .S0(n916[5]), .S1(n916[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_58_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_58_add_2_7.INJECT1_0 = "NO";
    defparam sub_58_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24282), 
          .COUT(n24283), .S0(n916[3]), .S1(n916[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_58_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_58_add_2_5.INJECT1_0 = "NO";
    defparam sub_58_add_2_5.INJECT1_1 = "NO";
    FD1P3AX valid_48 (.D(n27113), .SP(n24988), .CK(debug_c_c), .Q(n1009));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    CCU2D sub_58_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24281), 
          .COUT(n24282), .S0(n916[1]), .S1(n916[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_58_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_58_add_2_3.INJECT1_0 = "NO";
    defparam sub_58_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24281), 
          .S1(n916[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_58_add_2_1.INIT0 = 16'hF000;
    defparam sub_58_add_2_1.INIT1 = 16'h5555;
    defparam sub_58_add_2_1.INJECT1_0 = "NO";
    defparam sub_58_add_2_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U4
//

module PWMReceiver_U4 (GND_net, n27582, n27640, n28893, debug_c_c, 
            \register[2] , n12804, rc_ch2_c, n994, n24993) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n27582;
    output n27640;
    input n28893;
    input debug_c_c;
    output [7:0]\register[2] ;
    input n12804;
    input rc_ch2_c;
    output n994;
    input n24993;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n152, n103;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    
    wire n154, n24016, n29055;
    wire [15:0]n116;
    
    wire n24015, n29033, n24014, n29043, n24013, n29061, n29014, 
        n24012, n29060, n25137, n24992, n5, n27241, n27262, n27165, 
        n28993, n24851, n27021, n988, n1000, n27117, n24011, n28939, 
        n28967, n10, n11, n27315, n14411, n27018, n4, n4_adj_3, 
        n29062, n29013, n29064, n11790, n24010, n6;
    wire [7:0]n43;
    
    wire n24009, n28940, n27116, n4_adj_4, n28992;
    wire [7:0]n907;
    
    wire n24288, n24287, n24286, n24285;
    
    PFUMX i13582 (.BLUT(n152), .ALUT(n103), .C0(count[3]), .Z(n154));
    CCU2D add_1473_17 (.A0(count[15]), .B0(n29055), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24016), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_17.INIT0 = 16'hd222;
    defparam add_1473_17.INIT1 = 16'h0000;
    defparam add_1473_17.INJECT1_0 = "NO";
    defparam add_1473_17.INJECT1_1 = "NO";
    CCU2D add_1473_15 (.A0(count[13]), .B0(n29055), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n29055), .C1(GND_net), .D1(GND_net), .CIN(n24015), 
          .COUT(n24016), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_15.INIT0 = 16'hd222;
    defparam add_1473_15.INIT1 = 16'hd222;
    defparam add_1473_15.INJECT1_0 = "NO";
    defparam add_1473_15.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_375 (.A(count[7]), .B(count[6]), .C(count[8]), .Z(n29033)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_375.init = 16'hfefe;
    CCU2D add_1473_13 (.A0(count[11]), .B0(n29055), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n29055), .C1(GND_net), .D1(GND_net), .CIN(n24014), 
          .COUT(n24015), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_13.INIT0 = 16'hd222;
    defparam add_1473_13.INIT1 = 16'hd222;
    defparam add_1473_13.INJECT1_0 = "NO";
    defparam add_1473_13.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(count[7]), .B(count[6]), .C(count[8]), .D(n29043), 
         .Z(n103)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    CCU2D add_1473_11 (.A0(count[9]), .B0(n29055), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n29055), .C1(GND_net), .D1(GND_net), .CIN(n24013), 
          .COUT(n24014), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_11.INIT0 = 16'hd222;
    defparam add_1473_11.INIT1 = 16'hd222;
    defparam add_1473_11.INJECT1_0 = "NO";
    defparam add_1473_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_385 (.A(count[4]), .B(count[5]), .Z(n29043)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_rep_385.init = 16'h8888;
    LUT4 i1_3_lut_rep_356_4_lut (.A(count[4]), .B(count[5]), .C(n29061), 
         .D(count[3]), .Z(n29014)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_3_lut_rep_356_4_lut.init = 16'h8000;
    CCU2D add_1473_9 (.A0(count[7]), .B0(n29055), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n29055), .C1(GND_net), .D1(GND_net), .CIN(n24012), 
          .COUT(n24013), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_9.INIT0 = 16'hd222;
    defparam add_1473_9.INIT1 = 16'hd222;
    defparam add_1473_9.INJECT1_0 = "NO";
    defparam add_1473_9.INJECT1_1 = "NO";
    LUT4 i21299_4_lut (.A(n29060), .B(n29055), .C(n25137), .D(n24992), 
         .Z(n27582)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i21299_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n5), .B(n27241), .C(n27262), .D(n27165), .Z(n24992)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccec;
    LUT4 i20894_3_lut_4_lut (.A(count[8]), .B(n28993), .C(n24851), .D(n27021), 
         .Z(n27262)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i20894_3_lut_4_lut.init = 16'hfeee;
    LUT4 i5_2_lut_rep_397 (.A(n988), .B(n1000), .Z(n29055)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i5_2_lut_rep_397.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n988), .B(n1000), .C(n25137), .D(n29060), 
         .Z(n27117)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff4;
    CCU2D add_1473_7 (.A0(count[5]), .B0(n29055), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n29055), .C1(GND_net), .D1(GND_net), .CIN(n24011), 
          .COUT(n24012), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_7.INIT0 = 16'hd222;
    defparam add_1473_7.INIT1 = 16'hd222;
    defparam add_1473_7.INJECT1_0 = "NO";
    defparam add_1473_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_402 (.A(count[15]), .B(count[14]), .Z(n29060)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_402.init = 16'heeee;
    LUT4 i21357_4_lut (.A(n28939), .B(n27241), .C(n28967), .D(n10), 
         .Z(n27640)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i21357_4_lut.init = 16'h3323;
    LUT4 i2_4_lut (.A(n28893), .B(n29060), .C(n11), .D(n27315), .Z(n14411)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i2_4_lut.init = 16'h0020;
    LUT4 i4_4_lut (.A(n27018), .B(n27241), .C(n154), .D(count[9]), .Z(n11)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i4_4_lut.init = 16'h0322;
    LUT4 i1_2_lut_rep_403 (.A(count[2]), .B(count[1]), .Z(n29061)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_403.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[4]), .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[2]), .B(count[1]), .C(count[5]), .D(count[3]), 
         .Z(n4_adj_3)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_rep_404 (.A(count[7]), .B(count[6]), .Z(n29062)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_404.init = 16'h8888;
    LUT4 i1_2_lut_rep_355_3_lut (.A(count[7]), .B(count[6]), .C(count[8]), 
         .Z(n29013)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_355_3_lut.init = 16'h8080;
    LUT4 i20875_2_lut (.A(n988), .B(n1000), .Z(n27241)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i20875_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut_4_lut_adj_13 (.A(count[7]), .B(count[6]), .C(count[0]), 
         .D(n29014), .Z(n27021)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_3_lut_4_lut_adj_13.init = 16'h8000;
    LUT4 i2_4_lut_adj_14 (.A(n29062), .B(count[5]), .C(count[3]), .D(n4), 
         .Z(n24851)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_4_lut_adj_14.init = 16'h8880;
    LUT4 i3_4_lut (.A(count[12]), .B(count[13]), .C(n29060), .D(n29064), 
         .Z(n11790)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_406 (.A(count[10]), .B(count[11]), .Z(n29064)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_406.init = 16'heeee;
    LUT4 i20945_3_lut_4_lut (.A(count[10]), .B(count[11]), .C(count[13]), 
         .D(count[12]), .Z(n27315)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20945_3_lut_4_lut.init = 16'hfffe;
    LUT4 i20801_3_lut (.A(n11790), .B(count[9]), .C(n154), .Z(n27165)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i20801_3_lut.init = 16'heaea;
    CCU2D add_1473_5 (.A0(count[3]), .B0(n29055), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n29055), .C1(GND_net), .D1(GND_net), .CIN(n24010), 
          .COUT(n24011), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_5.INIT0 = 16'hd222;
    defparam add_1473_5.INIT1 = 16'hd222;
    defparam add_1473_5.INJECT1_0 = "NO";
    defparam add_1473_5.INJECT1_1 = "NO";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    LUT4 i23_4_lut (.A(n29033), .B(count[2]), .C(n29043), .D(n6), .Z(n152)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'hfaea;
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    LUT4 i2_2_lut (.A(count[1]), .B(count[0]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n12804), .PD(n14411), .CK(debug_c_c), 
            .Q(\register[2] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n12804), .PD(n14411), .CK(debug_c_c), 
            .Q(\register[2] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n12804), .PD(n14411), .CK(debug_c_c), 
            .Q(\register[2] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n12804), .PD(n14411), .CK(debug_c_c), 
            .Q(\register[2] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n12804), .PD(n14411), .CK(debug_c_c), 
            .Q(\register[2] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n12804), .PD(n14411), .CK(debug_c_c), 
            .Q(\register[2] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    CCU2D add_1473_3 (.A0(count[1]), .B0(n29055), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n29055), .C1(GND_net), .D1(GND_net), .CIN(n24009), 
          .COUT(n24010), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_3.INIT0 = 16'hd222;
    defparam add_1473_3.INIT1 = 16'hd222;
    defparam add_1473_3.INJECT1_0 = "NO";
    defparam add_1473_3.INJECT1_1 = "NO";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n12804), .PD(n14411), .CK(debug_c_c), 
            .Q(\register[2] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i21279_3_lut_3_lut_4_lut (.A(n29060), .B(n25137), .C(n28940), 
         .D(n27165), .Z(n27116)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i21279_3_lut_3_lut_4_lut.init = 16'h0010;
    IFS1P3DX latched_in_45 (.D(rc_ch2_c), .SP(n28893), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1000));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_15 (.A(count[13]), .B(count[12]), .C(n29064), .D(n4_adj_4), 
         .Z(n25137)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_15.init = 16'h8880;
    LUT4 i1_4_lut_adj_16 (.A(count[9]), .B(count[4]), .C(n29013), .D(n4_adj_3), 
         .Z(n4_adj_4)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_16.init = 16'hfaea;
    LUT4 i1_3_lut_rep_309_4_lut (.A(n29062), .B(n29014), .C(count[8]), 
         .D(n28993), .Z(n28967)) /* synthesis lut_function=(A (B+((D)+!C))+!A ((D)+!C)) */ ;
    defparam i1_3_lut_rep_309_4_lut.init = 16'hff8f;
    LUT4 i1_2_lut_rep_335 (.A(count[9]), .B(n11790), .Z(n28993)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i1_2_lut_rep_335.init = 16'heeee;
    LUT4 i21_3_lut_rep_281_4_lut (.A(count[9]), .B(n11790), .C(n27165), 
         .D(n27018), .Z(n28939)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i21_3_lut_rep_281_4_lut.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_282_3_lut_4_lut (.A(count[9]), .B(n11790), .C(n24851), 
         .D(count[8]), .Z(n28940)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i1_2_lut_rep_282_3_lut_4_lut.init = 16'hfffe;
    CCU2D add_1473_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n27117), .B1(n1000), .C1(count[0]), .D1(n988), .COUT(n24009), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_1.INIT0 = 16'hF000;
    defparam add_1473_1.INIT1 = 16'ha565;
    defparam add_1473_1.INJECT1_0 = "NO";
    defparam add_1473_1.INJECT1_1 = "NO";
    LUT4 i14536_2_lut_4_lut (.A(n28993), .B(count[8]), .C(n28992), .D(n907[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14536_2_lut_4_lut.init = 16'h0400;
    LUT4 i14535_2_lut_4_lut (.A(n28993), .B(count[8]), .C(n28992), .D(n907[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14535_2_lut_4_lut.init = 16'h0400;
    LUT4 i2_3_lut_4_lut (.A(count[8]), .B(n29062), .C(n29014), .D(count[0]), 
         .Z(n27018)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_3_lut_4_lut.init = 16'h8000;
    LUT4 i14534_2_lut_4_lut (.A(n28993), .B(count[8]), .C(n28992), .D(n907[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14534_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_rep_334_4_lut (.A(count[3]), .B(n29061), .C(n29043), 
         .D(n29062), .Z(n28992)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_rep_334_4_lut.init = 16'h8000;
    LUT4 i14533_2_lut_4_lut (.A(n28993), .B(count[8]), .C(n28992), .D(n907[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14533_2_lut_4_lut.init = 16'h0400;
    FD1P3AX prev_in_46 (.D(n1000), .SP(n28893), .CK(debug_c_c), .Q(n988));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut_adj_17 (.A(n27018), .B(n27165), .C(n28993), .D(n28967), 
         .Z(n5)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B !(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[13:39])
    defparam i1_2_lut_4_lut_adj_17.init = 16'hcd00;
    LUT4 i14532_2_lut_4_lut (.A(n28993), .B(count[8]), .C(n28992), .D(n907[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14532_2_lut_4_lut.init = 16'h0400;
    LUT4 i14531_2_lut_4_lut (.A(n28993), .B(count[8]), .C(n28992), .D(n907[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14531_2_lut_4_lut.init = 16'h0400;
    CCU2D sub_57_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24288), 
          .S0(n907[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_57_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_9.INIT1 = 16'h0000;
    defparam sub_57_add_2_9.INJECT1_0 = "NO";
    defparam sub_57_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24287), 
          .COUT(n24288), .S0(n907[5]), .S1(n907[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_57_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_57_add_2_7.INJECT1_0 = "NO";
    defparam sub_57_add_2_7.INJECT1_1 = "NO";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n12804), .PD(n14411), .CK(debug_c_c), 
            .Q(\register[2] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    CCU2D sub_57_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24286), 
          .COUT(n24287), .S0(n907[3]), .S1(n907[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_57_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_57_add_2_5.INJECT1_0 = "NO";
    defparam sub_57_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24285), 
          .COUT(n24286), .S0(n907[1]), .S1(n907[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_57_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_57_add_2_3.INJECT1_0 = "NO";
    defparam sub_57_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24285), 
          .S1(n907[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_57_add_2_1.INIT0 = 16'hF000;
    defparam sub_57_add_2_1.INIT1 = 16'h5555;
    defparam sub_57_add_2_1.INJECT1_0 = "NO";
    defparam sub_57_add_2_1.INJECT1_1 = "NO";
    LUT4 i14530_2_lut_4_lut (.A(n28993), .B(count[8]), .C(n28992), .D(n907[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14530_2_lut_4_lut.init = 16'h0400;
    FD1P3AX valid_48 (.D(n27116), .SP(n24993), .CK(debug_c_c), .Q(n994));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i14342_2_lut_4_lut (.A(n28993), .B(count[8]), .C(n28992), .D(n907[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14342_2_lut_4_lut.init = 16'h0400;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n28993), .C(n27021), 
         .D(n24851), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    
endmodule
//
// Verilog Description of module PWMReceiver_U5
//

module PWMReceiver_U5 (n27493, n27638, debug_c_c, n28893, GND_net, 
            \register[1] , n12807, rc_ch1_c, n979, n24976) /* synthesis syn_module_defined=1 */ ;
    output n27493;
    output n27638;
    input debug_c_c;
    input n28893;
    input GND_net;
    output [7:0]\register[1] ;
    input n12807;
    input rc_ch1_c;
    output n979;
    input n24976;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    
    wire n28994, n110, n23, n28942, n28941, n20591, n24866, n11798, 
        n27091, n11749, n112, n116, n4, n24846, n5, n6, n27191, 
        n25023, n29067, n27056, n29065, n28969, n29066, n28970, 
        n27219, n28995;
    wire [7:0]n898;
    wire [7:0]n43;
    
    wire n4_adj_1, n27093, n4_adj_2, n973, n985, n27119;
    wire [15:0]n1;
    
    wire n14414, n28971, n26731, n24292, n24291, n24290, n24289, 
        n27120, n24024, n24023, n24022, n24021, n24020, n24019, 
        n24018, n24017;
    
    LUT4 i1_4_lut (.A(count[8]), .B(n28994), .C(count[1]), .D(n110), 
         .Z(n23)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0222;
    LUT4 i2_4_lut (.A(n28942), .B(n23), .C(n28941), .D(n20591), .Z(n24866)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i2_4_lut.init = 16'heefe;
    LUT4 i3_4_lut (.A(count[12]), .B(count[13]), .C(n11798), .D(n27091), 
         .Z(n11749)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(count[15]), .B(count[14]), .Z(n11798)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_1 (.A(count[11]), .B(count[10]), .Z(n27091)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_1.init = 16'heeee;
    LUT4 i2_4_lut_adj_2 (.A(n112), .B(n116), .C(n4), .D(count[5]), .Z(n24846)) /* synthesis lut_function=(A (B (D))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i2_4_lut_adj_2.init = 16'hc800;
    LUT4 i1_2_lut_adj_3 (.A(count[4]), .B(count[3]), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_3.init = 16'heeee;
    LUT4 i20827_4_lut (.A(n11749), .B(count[9]), .C(n5), .D(n6), .Z(n27191)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i20827_4_lut.init = 16'heeea;
    LUT4 i2_2_lut (.A(count[6]), .B(count[8]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_4 (.A(count[0]), .B(count[3]), .C(count[1]), .D(count[2]), 
         .Z(n25023)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_4.init = 16'hfffe;
    LUT4 i1_2_lut_adj_5 (.A(count[2]), .B(count[1]), .Z(n112)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_5.init = 16'h8888;
    LUT4 i1_2_lut_adj_6 (.A(count[7]), .B(count[6]), .Z(n116)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_adj_6.init = 16'h8888;
    LUT4 i3_4_lut_adj_7 (.A(count[3]), .B(n116), .C(count[2]), .D(n29067), 
         .Z(n110)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i3_4_lut_adj_7.init = 16'h8000;
    LUT4 i21210_4_lut (.A(n27056), .B(n29065), .C(n28969), .D(n29066), 
         .Z(n27493)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i21210_4_lut.init = 16'h3031;
    LUT4 i4_4_lut (.A(n28970), .B(n27219), .C(n28995), .D(n24846), .Z(n27056)) /* synthesis lut_function=(!(A (B)+!A (B+!(C (D))))) */ ;
    defparam i4_4_lut.init = 16'h3222;
    LUT4 i14526_2_lut (.A(n898[6]), .B(n23), .Z(n43[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14526_2_lut.init = 16'h8888;
    LUT4 i14525_2_lut (.A(n898[5]), .B(n23), .Z(n43[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14525_2_lut.init = 16'h8888;
    LUT4 i14524_2_lut (.A(n898[4]), .B(n23), .Z(n43[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14524_2_lut.init = 16'h8888;
    LUT4 i14523_2_lut (.A(n898[3]), .B(n23), .Z(n43[3])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14523_2_lut.init = 16'h8888;
    LUT4 i14522_2_lut (.A(n898[2]), .B(n23), .Z(n43[2])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14522_2_lut.init = 16'h8888;
    LUT4 i14521_2_lut (.A(n898[1]), .B(n23), .Z(n43[1])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14521_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_8 (.A(n27091), .B(count[9]), .C(count[8]), .D(n4_adj_1), 
         .Z(n27093)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_8.init = 16'hfeee;
    LUT4 i1_4_lut_adj_9 (.A(n116), .B(count[3]), .C(n4_adj_2), .D(n112), 
         .Z(n4_adj_1)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_4_lut_adj_9.init = 16'ha8a0;
    LUT4 i1_2_lut_adj_10 (.A(count[4]), .B(count[5]), .Z(n4_adj_2)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_10.init = 16'heeee;
    LUT4 i5_2_lut_rep_407 (.A(n973), .B(n985), .Z(n29065)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i5_2_lut_rep_407.init = 16'h4444;
    LUT4 i1_2_lut_3_lut (.A(n973), .B(n985), .C(n28969), .Z(n27119)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i1_2_lut_3_lut.init = 16'hf4f4;
    LUT4 i1_2_lut_rep_408 (.A(n985), .B(n973), .Z(n29066)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_408.init = 16'hbbbb;
    LUT4 i21355_2_lut_3_lut (.A(n985), .B(n973), .C(n24866), .Z(n27638)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i21355_2_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_409 (.A(count[4]), .B(count[5]), .Z(n29067)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_rep_409.init = 16'h8888;
    LUT4 i1_3_lut_4_lut (.A(count[4]), .B(count[5]), .C(count[7]), .D(n25023), 
         .Z(n5)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    FD1P3IX count_i0_i15 (.D(n1[15]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n1[14]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n1[13]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n1[12]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n1[11]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n1[10]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n1[9]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n1[8]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n1[7]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n1[6]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n1[5]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n1[4]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n1[3]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n1[2]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n1[1]), .SP(n28893), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n12807), .PD(n14414), .CK(debug_c_c), 
            .Q(\register[1] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n12807), .PD(n14414), .CK(debug_c_c), 
            .Q(\register[1] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n12807), .PD(n14414), .CK(debug_c_c), 
            .Q(\register[1] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n12807), .PD(n14414), .CK(debug_c_c), 
            .Q(\register[1] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n12807), .PD(n14414), .CK(debug_c_c), 
            .Q(\register[1] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n12807), .PD(n14414), .CK(debug_c_c), 
            .Q(\register[1] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n12807), .PD(n14414), .CK(debug_c_c), 
            .Q(\register[1] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_336 (.A(count[9]), .B(n11749), .Z(n28994)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i1_2_lut_rep_336.init = 16'heeee;
    LUT4 i14846_2_lut_3_lut_4_lut (.A(count[9]), .B(n11749), .C(n28995), 
         .D(count[8]), .Z(n20591)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i14846_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_312_3_lut (.A(count[9]), .B(n11749), .C(count[8]), 
         .Z(n28970)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i1_2_lut_rep_312_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_283_3_lut_4_lut (.A(count[9]), .B(n11749), .C(n24846), 
         .D(count[8]), .Z(n28941)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i1_2_lut_rep_283_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_337 (.A(n110), .B(count[1]), .C(count[0]), .Z(n28995)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i2_3_lut_rep_337.init = 16'h8080;
    LUT4 i1_2_lut_rep_313_4_lut (.A(n110), .B(count[1]), .C(count[0]), 
         .D(count[8]), .Z(n28971)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_313_4_lut.init = 16'h8000;
    LUT4 i21_3_lut_rep_284_4_lut (.A(count[8]), .B(n28995), .C(n28994), 
         .D(n27191), .Z(n28942)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i21_3_lut_rep_284_4_lut.init = 16'h00f8;
    FD1P3AX prev_in_46 (.D(n985), .SP(n28893), .CK(debug_c_c), .Q(n973));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch1_c), .SP(n28893), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n985));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i3_4_lut_adj_11 (.A(n973), .B(n28893), .C(n26731), .D(n27191), 
         .Z(n14414)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut_adj_11.init = 16'h0080;
    LUT4 i2_4_lut_adj_12 (.A(n28971), .B(n24866), .C(count[9]), .D(n985), 
         .Z(n26731)) /* synthesis lut_function=(!(A ((D)+!B)+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i2_4_lut_adj_12.init = 16'h00c8;
    LUT4 i14336_2_lut (.A(n898[0]), .B(n23), .Z(n43[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14336_2_lut.init = 16'h8888;
    CCU2D sub_56_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24292), 
          .S0(n898[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_56_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_9.INIT1 = 16'h0000;
    defparam sub_56_add_2_9.INJECT1_0 = "NO";
    defparam sub_56_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_56_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24291), 
          .COUT(n24292), .S0(n898[5]), .S1(n898[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_56_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_56_add_2_7.INJECT1_0 = "NO";
    defparam sub_56_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_56_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24290), 
          .COUT(n24291), .S0(n898[3]), .S1(n898[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_56_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_56_add_2_5.INJECT1_0 = "NO";
    defparam sub_56_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_56_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24289), 
          .COUT(n24290), .S0(n898[1]), .S1(n898[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_56_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_56_add_2_3.INJECT1_0 = "NO";
    defparam sub_56_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_56_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24289), 
          .S1(n898[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_56_add_2_1.INIT0 = 16'hF000;
    defparam sub_56_add_2_1.INIT1 = 16'h5555;
    defparam sub_56_add_2_1.INJECT1_0 = "NO";
    defparam sub_56_add_2_1.INJECT1_1 = "NO";
    FD1P3IX count_i0_i0 (.D(n1[0]), .SP(n28893), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n12807), .PD(n14414), .CK(debug_c_c), 
            .Q(\register[1] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i14527_2_lut (.A(n898[7]), .B(n23), .Z(n43[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14527_2_lut.init = 16'h8888;
    FD1P3AX valid_48 (.D(n27120), .SP(n24976), .CK(debug_c_c), .Q(n979));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i21233_3_lut_3_lut_4_lut (.A(n24846), .B(n28970), .C(n27191), 
         .D(n28969), .Z(n27120)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i21233_3_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i20873_4_lut_rep_311 (.A(n11798), .B(count[13]), .C(count[12]), 
         .D(n27093), .Z(n28969)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i20873_4_lut_rep_311.init = 16'heaaa;
    CCU2D add_1469_17 (.A0(count[15]), .B0(n29065), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24024), 
          .S0(n1[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1469_17.INIT0 = 16'hd222;
    defparam add_1469_17.INIT1 = 16'h0000;
    defparam add_1469_17.INJECT1_0 = "NO";
    defparam add_1469_17.INJECT1_1 = "NO";
    CCU2D add_1469_15 (.A0(count[13]), .B0(n29065), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n29065), .C1(GND_net), .D1(GND_net), .CIN(n24023), 
          .COUT(n24024), .S0(n1[13]), .S1(n1[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1469_15.INIT0 = 16'hd222;
    defparam add_1469_15.INIT1 = 16'hd222;
    defparam add_1469_15.INJECT1_0 = "NO";
    defparam add_1469_15.INJECT1_1 = "NO";
    CCU2D add_1469_13 (.A0(count[11]), .B0(n29065), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n29065), .C1(GND_net), .D1(GND_net), .CIN(n24022), 
          .COUT(n24023), .S0(n1[11]), .S1(n1[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1469_13.INIT0 = 16'hd222;
    defparam add_1469_13.INIT1 = 16'hd222;
    defparam add_1469_13.INJECT1_0 = "NO";
    defparam add_1469_13.INJECT1_1 = "NO";
    CCU2D add_1469_11 (.A0(count[9]), .B0(n29065), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n29065), .C1(GND_net), .D1(GND_net), .CIN(n24021), 
          .COUT(n24022), .S0(n1[9]), .S1(n1[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1469_11.INIT0 = 16'hd222;
    defparam add_1469_11.INIT1 = 16'hd222;
    defparam add_1469_11.INJECT1_0 = "NO";
    defparam add_1469_11.INJECT1_1 = "NO";
    CCU2D add_1469_9 (.A0(count[7]), .B0(n29065), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n29065), .C1(GND_net), .D1(GND_net), .CIN(n24020), 
          .COUT(n24021), .S0(n1[7]), .S1(n1[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1469_9.INIT0 = 16'hd222;
    defparam add_1469_9.INIT1 = 16'hd222;
    defparam add_1469_9.INJECT1_0 = "NO";
    defparam add_1469_9.INJECT1_1 = "NO";
    CCU2D add_1469_7 (.A0(count[5]), .B0(n29065), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n29065), .C1(GND_net), .D1(GND_net), .CIN(n24019), 
          .COUT(n24020), .S0(n1[5]), .S1(n1[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1469_7.INIT0 = 16'hd222;
    defparam add_1469_7.INIT1 = 16'hd222;
    defparam add_1469_7.INJECT1_0 = "NO";
    defparam add_1469_7.INJECT1_1 = "NO";
    CCU2D add_1469_5 (.A0(count[3]), .B0(n29065), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n29065), .C1(GND_net), .D1(GND_net), .CIN(n24018), 
          .COUT(n24019), .S0(n1[3]), .S1(n1[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1469_5.INIT0 = 16'hd222;
    defparam add_1469_5.INIT1 = 16'hd222;
    defparam add_1469_5.INJECT1_0 = "NO";
    defparam add_1469_5.INJECT1_1 = "NO";
    LUT4 i20854_3_lut_4_lut (.A(n28971), .B(n27191), .C(n28994), .D(n23), 
         .Z(n27219)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[13:39])
    defparam i20854_3_lut_4_lut.init = 16'hfffe;
    CCU2D add_1469_3 (.A0(count[1]), .B0(n29065), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n29065), .C1(GND_net), .D1(GND_net), .CIN(n24017), 
          .COUT(n24018), .S0(n1[1]), .S1(n1[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1469_3.INIT0 = 16'hd222;
    defparam add_1469_3.INIT1 = 16'hd222;
    defparam add_1469_3.INJECT1_0 = "NO";
    defparam add_1469_3.INJECT1_1 = "NO";
    CCU2D add_1469_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n27119), .B1(n985), .C1(count[0]), .D1(n973), .COUT(n24017), 
          .S1(n1[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1469_1.INIT0 = 16'hF000;
    defparam add_1469_1.INIT1 = 16'ha565;
    defparam add_1469_1.INJECT1_0 = "NO";
    defparam add_1469_1.INJECT1_1 = "NO";
    
endmodule

// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.4.1.213
// Netlist written on Mon Jan 18 16:24:47 2016
//
// Verilog Description of module UniboardTop
//

module UniboardTop (uart_rx, uart_tx, status_led, clk_12MHz, Stepper_X_Step, 
            Stepper_X_Dir, Stepper_X_M0, Stepper_X_M1, Stepper_X_M2, 
            Stepper_X_En, Stepper_X_nFault, Stepper_Y_Step, Stepper_Y_Dir, 
            Stepper_Y_M0, Stepper_Y_M1, Stepper_Y_M2, Stepper_Y_En, 
            Stepper_Y_nFault, Stepper_Z_Step, Stepper_Z_Dir, Stepper_Z_M0, 
            Stepper_Z_M1, Stepper_Z_M2, Stepper_Z_En, Stepper_Z_nFault, 
            Stepper_A_Step, Stepper_A_Dir, Stepper_A_M0, Stepper_A_M1, 
            Stepper_A_M2, Stepper_A_En, Stepper_A_nFault, limit, expansion1, 
            expansion2, expansion3, expansion4, expansion5, signal_light, 
            encoder_ra, encoder_rb, encoder_ri, encoder_la, encoder_lb, 
            encoder_li, rc_ch1, rc_ch2, rc_ch3, rc_ch4, rc_ch7, 
            rc_ch8, motor_pwm_l, motor_pwm_r, xbee_pause, debug) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(363[8:19])
    input uart_rx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[13:20])
    output uart_tx;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[14:21])
    output [2:0]status_led;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    input clk_12MHz;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    output Stepper_X_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:31])
    output Stepper_X_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:30])
    output Stepper_X_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    output Stepper_X_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    output Stepper_X_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    output Stepper_X_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[17:29])
    input Stepper_X_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(375[16:32])
    output Stepper_Y_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:31])
    output Stepper_Y_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:30])
    output Stepper_Y_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    output Stepper_Y_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    output Stepper_Y_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    output Stepper_Y_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[17:29])
    input Stepper_Y_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(383[16:32])
    output Stepper_Z_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:31])
    output Stepper_Z_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:30])
    output Stepper_Z_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    output Stepper_Z_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    output Stepper_Z_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    output Stepper_Z_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[17:29])
    input Stepper_Z_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(391[16:32])
    output Stepper_A_Step;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:31])
    output Stepper_A_Dir;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:30])
    output Stepper_A_M0;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    output Stepper_A_M1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    output Stepper_A_M2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    output Stepper_A_En;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[17:29])
    input Stepper_A_nFault;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(399[16:32])
    input [3:0]limit;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    output expansion1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    output expansion2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    output expansion3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[14:24])
    output expansion4 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    output expansion5 /* synthesis .original_dir=IN_OUT */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[13:23])
    output signal_light;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(407[14:26])
    input encoder_ra;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(409[13:23])
    input encoder_rb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(410[13:23])
    input encoder_ri;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(411[13:23])
    input encoder_la;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(412[13:23])
    input encoder_lb;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(413[13:23])
    input encoder_li;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(414[13:23])
    input rc_ch1;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    input rc_ch2;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    input rc_ch3;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    input rc_ch4;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    input rc_ch7;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    input rc_ch8;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(421[13:19])
    output motor_pwm_l;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    output motor_pwm_r;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[14:25])
    input xbee_pause;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(425[13:23])
    output [8:0]debug;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [127:0]select /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    
    wire GND_net, VCC_net, n9396_c, n9395, Stepper_X_Step_c, Stepper_X_Dir_c, 
        Stepper_X_M0_c_0, Stepper_X_M1_c_1, Stepper_X_M2_c_2, Stepper_X_En_c, 
        Stepper_X_nFault_c, Stepper_Y_Step_c, Stepper_Y_Dir_c, Stepper_Y_M0_c_0, 
        Stepper_Y_M1_c_1, Stepper_Y_M2_c_2, Stepper_Y_En_c, Stepper_Y_nFault_c, 
        Stepper_Z_Step_c, Stepper_Z_Dir_c, Stepper_Z_M0_c_0, Stepper_Z_M1_c_1, 
        Stepper_Z_M2_c_2, Stepper_Z_En_c, Stepper_Z_nFault_c, Stepper_A_Step_c, 
        Stepper_A_Dir_c, Stepper_A_M0_c_0, Stepper_A_M1_c_1, Stepper_A_M2_c_2, 
        Stepper_A_En_c, Stepper_A_nFault_c, limit_c_3, limit_c_2, limit_c_1, 
        limit_c_0, signal_light_c, rc_ch1_c, rc_ch2_c, rc_ch3_c, rc_ch4_c, 
        rc_ch7_c, rc_ch8_c, xbee_pause_c, debug_c_7, debug_c_5, debug_c_4, 
        debug_c_3, debug_c_2;
    wire [31:0]databus;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(458[14:21])
    wire [2:0]reg_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(459[13:21])
    wire [7:0]register_addr;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    
    wire rw, n17, n15, n28324, n18770, n14, n15_adj_395;
    wire [15:0]reset_count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(465[13:24])
    wire [4:0]arm_select;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(524[12:22])
    
    wire n14473, n32371, n20505, n28332, n12620, n12434, n6, n29618, 
        n6_adj_396, n14446, n31426, n21, n10513, n31000, n1;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    wire [31:0]databus_out;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(55[13:24])
    
    wire n27764, n4, n27763, n2, n27762, n27761, n32369, n27760, 
        n27759;
    wire [31:0]n1286;
    
    wire n29663, n27758, n28304, n30866, n183, n2_adj_397, n28296, 
        n11753, n32366, n32365, force_pause;
    wire [31:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    wire [31:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    wire [31:0]read_value;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(30[13:23])
    wire [2:0]read_size;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(31[12:21])
    
    wire n12224;
    wire [7:0]n7893;
    
    wire n13, n11645, n1_adj_398, n2_adj_399, n30905, n9633, n30, 
        n15_adj_400, n241;
    wire [7:0]read_value_adj_690;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(63[12:22])
    wire [2:0]read_size_adj_691;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(64[12:21])
    
    wire n64;
    wire [15:0]n281;
    
    wire n30458;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    wire [31:0]read_value_adj_695;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_696;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select, n3363;
    wire [31:0]n224;
    
    wire n2_adj_444, n302;
    wire [31:0]n3451;
    
    wire n30338;
    wire [7:0]n571;
    
    wire n14322;
    wire [31:0]n580;
    
    wire n12138;
    wire [7:0]control_reg_adj_704;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]steps_reg_adj_706;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire stepping;
    wire [31:0]read_value_adj_707;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_708;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire n52, n32360, n7912, n32358, n32357, n32356, n19877, n30456;
    wire [7:0]control_reg_adj_744;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]steps_reg_adj_746;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire stepping_adj_483;
    wire [31:0]read_value_adj_747;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_748;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_518, n32354, n30995, n32353, n30969, n30284;
    wire [31:0]n3181;
    
    wire n3589, n32352, n12098, n16, motor_pwm_l_c, n4_adj_519, 
        n1_adj_520;
    wire [7:0]control_reg_adj_784;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [31:0]div_factor_reg_adj_785;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg_adj_786;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire stepping_adj_524;
    wire [31:0]read_value_adj_787;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(50[13:23])
    wire [2:0]read_size_adj_788;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(51[12:21])
    
    wire prev_select_adj_559, n3586;
    wire [31:0]n224_adj_791;
    
    wire n32350, n14_adj_592, n12, n2_adj_593, n27962, n10, n31427, 
        n32348, n28270, n12031, n12030, bclk;
    wire [7:0]rdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(22[12:17])
    wire [5:0]state_adj_834;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    
    wire n7852, n30310, n6_adj_594, n34317, n31049, n30240, n30710, 
        n4_adj_595, n32336, n6_adj_596, n5, n15_adj_597, n30911, 
        n30868, n32513, n4_adj_598, n28309, n34326, n28317, n30867, 
        n11981, n11966, n28312, n15_adj_599, n21_adj_600, n32505, 
        n32504, n32503, n2_adj_601, n30726, n30631, n4_adj_602, 
        n32495, n32494, n2_adj_603, n1_adj_604, n4_adj_605, n32486;
    wire [14:0]n66_adj_1129;
    
    wire n4_adj_606, n4_adj_607, n1_adj_608, n6_adj_609, n16_adj_610, 
        n14_adj_611, n12_adj_612, n10_adj_613, n8, n6_adj_614, n5_adj_615, 
        n4_adj_616, n32481, n4_adj_617, n32480, n4_adj_618, n1_adj_619, 
        n2_adj_620, n1_adj_621, n2_adj_622, n1_adj_623, n2_adj_624, 
        n1_adj_625, n2_adj_626, n34325, n32472, n4_adj_627, n1_adj_628, 
        n2_adj_629, n1_adj_630, n2_adj_631, n1_adj_632, n2_adj_633, 
        n1_adj_634, n2_adj_635, n1_adj_636, n2_adj_637, n32460, n1_adj_638, 
        n2_adj_639, n1_adj_640, n2_adj_641, n34324, n32455, n1_adj_642, 
        n2_adj_643, n1_adj_644, n2_adj_645, n1_adj_646, n32454, n30401, 
        n34323, n6_adj_647, n5_adj_648, n29158, n28308, n1_adj_649;
    wire [31:0]n6096;
    
    wire n32448, n32444, n14_adj_650, n32443, n2_adj_651, n32442, 
        n1_adj_652, n34322, n32440, n32439, n1_adj_653, n28459;
    wire [12:0]count_adj_845;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    
    wire n20268, n32345;
    wire [12:0]count_adj_848;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    wire [7:0]n7903;
    
    wire motor_pwm_r_c, n8_adj_661, n32433, n32432, n11883, n32429, 
        n31005, n32343, n30457, n32, n34321, n30913, n30810, n1_adj_662, 
        n2_adj_663, n32422, n30427, n30423, n30411, n7902, n32417, 
        n30802, n31442, n31441, n30797, n12841, n2_adj_664, n32412, 
        n32411, n30313, n32410, n30283, n32409, n32408, n8048, 
        n30929, n28356, n34320, n30258, n30211, n54, n20395, n32401, 
        n32399, n14_adj_665, n32398, n30787, n12788, n1_adj_666, 
        n2_adj_667, n1_adj_668, n30779, n32390, n32389, n6674, n32384, 
        n15_adj_669, n32383, n30774, n31024, n32381, n9, n32379, 
        n32341, n32376, n32375, n32374, n988, n32373, n1000, n11271;
    
    VHI i2 (.Z(VCC_net));
    PWMPeripheral motor_pwm (.\read_size[0] (read_size_adj_691[0]), .debug_c_c(debug_c_c), 
            .n30726(n30726), .n34322(n34322), .\databus[0] (databus[0]), 
            .\select[2] (select[2]), .rw(rw), .n32440(n32440), .\register_addr[0] (register_addr[0]), 
            .read_value({read_value_adj_690}), .n282(n281[15]), .n34326(n34326), 
            .\databus[6] (databus[6]), .\databus[5] (databus[5]), .\databus[4] (databus[4]), 
            .\databus[3] (databus[3]), .\databus[2] (databus[2]), .\databus[1] (databus[1]), 
            .n32448(n32448), .n32460(n32460), .n34320(n34320), .n34317(n34317), 
            .n64(n64), .\count[0] (count_adj_848[0]), .n32341(n32341), 
            .motor_pwm_r_c(motor_pwm_r_c), .GND_net(GND_net), .n9633(n9633), 
            .n14322(n14322), .\count[1] (count_adj_848[1]), .\count[2] (count_adj_848[2]), 
            .\count[3] (count_adj_848[3]), .\count[4] (count_adj_848[4]), 
            .\count[5] (count_adj_848[5]), .\count[6] (count_adj_848[6]), 
            .\count[7] (count_adj_848[7]), .\count[8] (count_adj_848[8]), 
            .n3589(n3589), .n7893({n7893}), .n7902(n7902), .n10513(n10513), 
            .n14473(n14473), .\count[0]_adj_195 (count_adj_845[0]), .\count[12] (count_adj_845[12]), 
            .\count[11] (count_adj_845[11]), .\count[9] (count_adj_845[9]), 
            .\count[8]_adj_196 (count_adj_845[8]), .\count[6]_adj_197 (count_adj_845[6]), 
            .\count[5]_adj_198 (count_adj_845[5]), .\count[3]_adj_199 (count_adj_845[3]), 
            .\count[2]_adj_200 (count_adj_845[2]), .\count[1]_adj_201 (count_adj_845[1]), 
            .motor_pwm_l_c(motor_pwm_l_c), .n28459(n28459), .n32356(n32356), 
            .n10(n10_adj_613), .n12(n12_adj_612), .\reset_count[6] (reset_count[6]), 
            .n30456(n30456), .\reset_count[4] (reset_count[4]), .\reset_count[5] (reset_count[5]), 
            .n30458(n30458), .\reset_count[12] (reset_count[12]), .\reset_count[11] (reset_count[11]), 
            .\reset_count[13] (reset_count[13]), .n29618(n29618), .n3586(n3586), 
            .n6(n6_adj_594), .n32411(n32411), .n6_adj_202(n6_adj_614), 
            .n8(n8), .n7912(n7912), .n7906(n7903[5]), .n7905(n7903[6]), 
            .n7908(n7903[3]), .n7910(n7903[1]), .n7909(n7903[2]), .n7911(n7903[0])) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(512[16] 522[40])
    LUT4 n227_bdd_4_lut (.A(n9396_c), .B(state_adj_834[1]), .C(rdata[0]), 
         .D(bclk), .Z(n31426)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C)+!B !((D)+!C))) */ ;
    defparam n227_bdd_4_lut.init = 16'he2f0;
    PFUMX i24509 (.BLUT(n30866), .ALUT(n30867), .C0(register_addr[1]), 
          .Z(n30868));
    PFUMX LessThan_1437_i18 (.BLUT(n14_adj_592), .ALUT(n16), .C0(n30810), 
          .Z(n3589));
    PFUMX LessThan_1434_i18 (.BLUT(n14_adj_611), .ALUT(n16_adj_610), .C0(n30787), 
          .Z(n3586));
    PFUMX i22 (.BLUT(n15_adj_597), .ALUT(n30905), .C0(state_adj_834[0]), 
          .Z(n29158));
    LUT4 i2_2_lut_rep_315_3_lut_4_lut (.A(n32495), .B(n32494), .C(state_adj_834[5]), 
         .D(state_adj_834[0]), .Z(n32409)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i2_2_lut_rep_315_3_lut_4_lut.init = 16'h0010;
    LUT4 LessThan_1434_i11_2_lut_rep_290 (.A(n7903[5]), .B(count_adj_845[5]), 
         .Z(n32384)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i11_2_lut_rep_290.init = 16'h6666;
    LUT4 i13936_2_lut_2_lut (.A(n34320), .B(n6674), .Z(n241)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i13936_2_lut_2_lut.init = 16'h4444;
    LUT4 LessThan_1437_i13_2_lut_rep_277 (.A(n7893[6]), .B(count_adj_848[6]), 
         .Z(n32371)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i13_2_lut_rep_277.init = 16'h6666;
    LUT4 LessThan_1437_i10_3_lut_3_lut (.A(n7893[6]), .B(count_adj_848[6]), 
         .C(count_adj_848[5]), .Z(n10)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i10_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i13975_2_lut_2_lut (.A(n34320), .B(databus[7]), .Z(n281[15])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i13975_2_lut_2_lut.init = 16'h4444;
    LUT4 LessThan_1437_i11_2_lut_rep_279 (.A(n7893[5]), .B(count_adj_848[5]), 
         .Z(n32373)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i11_2_lut_rep_279.init = 16'h6666;
    PFUMX i13028 (.BLUT(n18770), .ALUT(n15), .C0(register_addr[0]), .Z(n6096[4]));
    LUT4 i24443_2_lut_3_lut_4_lut (.A(n7893[5]), .B(count_adj_848[5]), .C(count_adj_848[6]), 
         .D(n7893[6]), .Z(n30802)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24443_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i13026_3_lut (.A(control_reg_adj_784[4]), .B(div_factor_reg_adj_785[4]), 
         .C(register_addr[1]), .Z(n18770)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13026_3_lut.init = 16'hcaca;
    LUT4 n32503_bdd_4_lut (.A(n32503), .B(n32504), .C(register_addr[1]), 
         .D(register_addr[0]), .Z(n30423)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam n32503_bdd_4_lut.init = 16'h0010;
    LUT4 i24695_4_lut_rep_425 (.A(reset_count[14]), .B(n30458), .C(n29618), 
         .D(n19877), .Z(n34320)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24695_4_lut_rep_425.init = 16'h575f;
    LUT4 i24695_4_lut_rep_426 (.A(reset_count[14]), .B(n30458), .C(n29618), 
         .D(n19877), .Z(n34321)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24695_4_lut_rep_426.init = 16'h575f;
    LUT4 i2_3_lut (.A(reset_count[7]), .B(reset_count[5]), .C(reset_count[6]), 
         .Z(n27962)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i24695_4_lut_rep_427 (.A(reset_count[14]), .B(n30458), .C(n29618), 
         .D(n19877), .Z(n34322)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24695_4_lut_rep_427.init = 16'h575f;
    LUT4 i24695_4_lut_rep_428 (.A(reset_count[14]), .B(n30458), .C(n29618), 
         .D(n19877), .Z(n34323)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24695_4_lut_rep_428.init = 16'h575f;
    LUT4 i24420_2_lut_3_lut_4_lut (.A(n7903[5]), .B(count_adj_845[5]), .C(count_adj_845[6]), 
         .D(n7903[6]), .Z(n30779)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24420_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 Select_3607_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[13]), 
         .D(rw), .Z(n2_adj_631)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3607_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3595_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[19]), 
         .D(rw), .Z(n1_adj_634)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3595_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3603_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[15]), 
         .D(rw), .Z(n1_adj_642)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3603_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3609_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[12]), 
         .D(rw), .Z(n2_adj_629)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3609_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3605_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[14]), 
         .D(rw), .Z(n1_adj_632)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3605_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i24695_4_lut_rep_429 (.A(reset_count[14]), .B(n30458), .C(n29618), 
         .D(n19877), .Z(n34324)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24695_4_lut_rep_429.init = 16'h575f;
    LUT4 i1_2_lut_rep_386 (.A(register_addr[4]), .B(register_addr[5]), .Z(n32480)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(527[4] 556[11])
    defparam i1_2_lut_rep_386.init = 16'heeee;
    FD1P3AX reset_count_2172_2173__i1 (.D(n66_adj_1129[0]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i1.GSR = "ENABLED";
    LUT4 Select_3607_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[13]), 
         .D(rw), .Z(n1_adj_630)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3607_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3609_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[12]), 
         .D(n34317), .Z(n1_adj_628)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3609_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_2_lut_rep_349_3_lut_4_lut (.A(register_addr[4]), .B(register_addr[5]), 
         .C(n32504), .D(n32481), .Z(n32443)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(527[4] 556[11])
    defparam i2_2_lut_rep_349_3_lut_4_lut.init = 16'hfffe;
    LUT4 i24236_2_lut_rep_335_3_lut_4_lut (.A(register_addr[4]), .B(register_addr[5]), 
         .C(register_addr[0]), .D(n32481), .Z(n32429)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(527[4] 556[11])
    defparam i24236_2_lut_rep_335_3_lut_4_lut.init = 16'hfffe;
    LUT4 Select_3611_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[11]), 
         .D(n34317), .Z(n1_adj_623)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3611_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3613_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[10]), 
         .D(n34317), .Z(n1_adj_619)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3613_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i24695_4_lut_rep_430 (.A(reset_count[14]), .B(n30458), .C(n29618), 
         .D(n19877), .Z(n34325)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24695_4_lut_rep_430.init = 16'h575f;
    LUT4 i1_4_lut (.A(div_factor_reg_adj_785[8]), .B(register_addr[1]), 
         .C(steps_reg_adj_786[8]), .D(register_addr[0]), .Z(n30211)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i24695_4_lut_rep_431 (.A(reset_count[14]), .B(n30458), .C(n29618), 
         .D(n19877), .Z(n34326)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24695_4_lut_rep_431.init = 16'h575f;
    LUT4 LessThan_1437_i15_2_lut_rep_258 (.A(n7893[7]), .B(count_adj_848[7]), 
         .Z(n32352)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i15_2_lut_rep_258.init = 16'h6666;
    LUT4 Select_3615_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[9]), 
         .D(rw), .Z(n1_adj_625)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3615_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 LessThan_1437_i12_3_lut_3_lut (.A(n7893[7]), .B(count_adj_848[7]), 
         .C(n10), .Z(n12)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i12_3_lut_3_lut.init = 16'hd4d4;
    LUT4 Select_3617_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[8]), 
         .D(rw), .Z(n1_adj_621)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3617_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 LessThan_1437_i17_2_lut_rep_259 (.A(n7902), .B(count_adj_848[8]), 
         .Z(n32353)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i17_2_lut_rep_259.init = 16'h6666;
    LUT4 Select_3611_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[11]), 
         .D(rw), .Z(n2_adj_624)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3611_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 LessThan_1437_i16_3_lut_3_lut (.A(n7902), .B(count_adj_848[8]), 
         .C(n8_adj_661), .Z(n16)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i16_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i24695_4_lut_rep_339 (.A(reset_count[14]), .B(n30458), .C(n29618), 
         .D(n19877), .Z(n32433)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C)))) */ ;
    defparam i24695_4_lut_rep_339.init = 16'h575f;
    LUT4 Select_3613_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[10]), 
         .D(rw), .Z(n2_adj_620)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3613_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 LessThan_1434_i17_2_lut_rep_263 (.A(n7912), .B(count_adj_845[8]), 
         .Z(n32357)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i17_2_lut_rep_263.init = 16'h6666;
    LUT4 Select_3615_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[9]), 
         .D(rw), .Z(n2_adj_626)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3615_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 LessThan_1434_i16_3_lut_3_lut (.A(n7912), .B(count_adj_845[8]), 
         .C(n8), .Z(n16_adj_610)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i16_3_lut_3_lut.init = 16'hd4d4;
    LUT4 Select_3571_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[31]), 
         .D(rw), .Z(n1_adj_604)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3571_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3617_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[8]), 
         .D(rw), .Z(n2_adj_622)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3617_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_rep_275_3_lut_4_lut (.A(n32454), .B(select[4]), .C(prev_select), 
         .D(n32480), .Z(n32369)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_275_3_lut_4_lut.init = 16'h0004;
    LUT4 i20_2_lut_rep_281_3_lut_4_lut (.A(n32454), .B(select[4]), .C(n34317), 
         .D(n32480), .Z(n32375)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i20_2_lut_rep_281_3_lut_4_lut.init = 16'h0040;
    LUT4 i20_2_lut_rep_280_3_lut_4_lut (.A(n32454), .B(select[4]), .C(rw), 
         .D(n30427), .Z(n32374)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i20_2_lut_rep_280_3_lut_4_lut.init = 16'h4000;
    LUT4 n9396_c_bdd_4_lut (.A(n9396_c), .B(state_adj_834[1]), .C(rdata[1]), 
         .D(bclk), .Z(n31441)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(B ((D)+!C)+!B !(C))) */ ;
    defparam n9396_c_bdd_4_lut.init = 16'hb8f0;
    LUT4 Select_3571_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[31]), 
         .D(rw), .Z(n2_adj_603)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3571_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i24806_4_lut (.A(n32357), .B(n32356), .C(n32383), .D(n30774), 
         .Z(n30787)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24806_4_lut.init = 16'habaa;
    LUT4 i1_2_lut_rep_287_3_lut_4_lut (.A(n32454), .B(select[4]), .C(prev_select_adj_559), 
         .D(n30427), .Z(n32381)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_rep_287_3_lut_4_lut.init = 16'h0400;
    LUT4 i20_2_lut_rep_282_3_lut_4_lut (.A(n32454), .B(select[4]), .C(rw), 
         .D(n32505), .Z(n32376)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i20_2_lut_rep_282_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_296_3_lut_4_lut (.A(n32454), .B(select[4]), .C(prev_select_adj_518), 
         .D(n32505), .Z(n32390)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_296_3_lut_4_lut.init = 16'h0004;
    LUT4 Select_3577_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[28]), 
         .D(rw), .Z(n1_adj_652)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3577_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_472 (.A(register_addr[1]), .B(div_factor_reg_adj_785[16]), 
         .C(steps_reg_adj_786[16]), .D(register_addr[0]), .Z(n17)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_472.init = 16'ha088;
    LUT4 i1_2_lut_rep_400 (.A(state_adj_834[1]), .B(state_adj_834[4]), .Z(n32494)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i1_2_lut_rep_400.init = 16'heeee;
    LUT4 i1_2_lut_rep_338_3_lut_4_lut (.A(state_adj_834[1]), .B(state_adj_834[4]), 
         .C(state_adj_834[0]), .D(n32495), .Z(n32432)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i1_2_lut_rep_338_3_lut_4_lut.init = 16'hfffe;
    LUT4 Select_3577_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[28]), 
         .D(rw), .Z(n2_adj_444)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3577_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state_adj_834[1]), .B(state_adj_834[4]), 
         .C(n9396_c), .D(n32495), .Z(n183)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_401 (.A(state_adj_834[2]), .B(state_adj_834[3]), .Z(n32495)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i1_2_lut_rep_401.init = 16'heeee;
    LUT4 Select_3573_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[30]), 
         .D(n34317), .Z(n1_adj_649)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3573_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 n31441_bdd_3_lut_4_lut (.A(state_adj_834[2]), .B(state_adj_834[3]), 
         .C(rdata[1]), .D(n31441), .Z(n31442)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam n31441_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n31426_bdd_3_lut_4_lut (.A(state_adj_834[2]), .B(state_adj_834[3]), 
         .C(rdata[0]), .D(n31426), .Z(n31427)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam n31426_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 Select_3575_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[29]), 
         .D(n34317), .Z(n1_adj_520)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3575_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3573_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[30]), 
         .D(rw), .Z(n2_adj_601)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3573_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3575_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[29]), 
         .D(rw), .Z(n2_adj_664)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3575_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    IB xbee_pause_pad (.I(xbee_pause), .O(xbee_pause_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(425[13:23])
    IB rc_ch8_pad (.I(rc_ch8), .O(rc_ch8_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(421[13:19])
    IB rc_ch7_pad (.I(rc_ch7), .O(rc_ch7_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(420[13:19])
    IB rc_ch4_pad (.I(rc_ch4), .O(rc_ch4_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(419[13:19])
    IB rc_ch3_pad (.I(rc_ch3), .O(rc_ch3_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(418[13:19])
    IB rc_ch2_pad (.I(rc_ch2), .O(rc_ch2_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(417[13:19])
    IB rc_ch1_pad (.I(rc_ch1), .O(rc_ch1_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(416[13:19])
    IB limit_pad_0 (.I(limit[0]), .O(limit_c_0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_1 (.I(limit[1]), .O(limit_c_1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_2 (.I(limit[2]), .O(limit_c_2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB limit_pad_3 (.I(limit[3]), .O(limit_c_3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(401[19:24])
    IB Stepper_A_nFault_pad (.I(Stepper_A_nFault), .O(Stepper_A_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(399[16:32])
    IB Stepper_Z_nFault_pad (.I(Stepper_Z_nFault), .O(Stepper_Z_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(391[16:32])
    IB Stepper_Y_nFault_pad (.I(Stepper_Y_nFault), .O(Stepper_Y_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(383[16:32])
    IB Stepper_X_nFault_pad (.I(Stepper_X_nFault), .O(Stepper_X_nFault_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(375[16:32])
    IB debug_c_pad (.I(clk_12MHz), .O(debug_c_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    IB n9396_pad (.I(uart_rx), .O(n9396_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(364[13:20])
    OB debug_pad_0 (.I(n9396_c), .O(debug[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_1 (.I(n9395), .O(debug[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_2 (.I(debug_c_2), .O(debug[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_3 (.I(debug_c_3), .O(debug[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_4 (.I(debug_c_4), .O(debug[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_5 (.I(debug_c_5), .O(debug[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_6 (.I(n34320), .O(debug[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_7 (.I(debug_c_7), .O(debug[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB debug_pad_8 (.I(debug_c_c), .O(debug[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(427[19:24])
    OB motor_pwm_r_pad (.I(motor_pwm_r_c), .O(motor_pwm_r));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(424[14:25])
    OB motor_pwm_l_pad (.I(motor_pwm_l_c), .O(motor_pwm_l));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(423[14:25])
    OB signal_light_pad (.I(signal_light_c), .O(signal_light));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(407[14:26])
    OB expansion5_pad (.I(GND_net), .O(expansion5));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(406[13:23])
    OB expansion4_pad (.I(GND_net), .O(expansion4));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(405[13:23])
    OB expansion3_pad (.I(GND_net), .O(expansion3));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(404[14:24])
    OB expansion2_pad (.I(GND_net), .O(expansion2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(403[14:24])
    OB expansion1_pad (.I(GND_net), .O(expansion1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(402[14:24])
    OB Stepper_A_En_pad (.I(Stepper_A_En_c), .O(Stepper_A_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(398[17:29])
    OB Stepper_A_M2_pad (.I(Stepper_A_M2_c_2), .O(Stepper_A_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(397[17:29])
    OB Stepper_A_M1_pad (.I(Stepper_A_M1_c_1), .O(Stepper_A_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(396[17:29])
    OB Stepper_A_M0_pad (.I(Stepper_A_M0_c_0), .O(Stepper_A_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(395[17:29])
    OB Stepper_A_Dir_pad (.I(Stepper_A_Dir_c), .O(Stepper_A_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(394[17:30])
    OB Stepper_A_Step_pad (.I(Stepper_A_Step_c), .O(Stepper_A_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(393[17:31])
    OB Stepper_Z_En_pad (.I(Stepper_Z_En_c), .O(Stepper_Z_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(390[17:29])
    OB Stepper_Z_M2_pad (.I(Stepper_Z_M2_c_2), .O(Stepper_Z_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(389[17:29])
    OB Stepper_Z_M1_pad (.I(Stepper_Z_M1_c_1), .O(Stepper_Z_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(388[17:29])
    OB Stepper_Z_M0_pad (.I(Stepper_Z_M0_c_0), .O(Stepper_Z_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(387[17:29])
    OB Stepper_Z_Dir_pad (.I(Stepper_Z_Dir_c), .O(Stepper_Z_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(386[17:30])
    OB Stepper_Z_Step_pad (.I(Stepper_Z_Step_c), .O(Stepper_Z_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(385[17:31])
    OB Stepper_Y_En_pad (.I(Stepper_Y_En_c), .O(Stepper_Y_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(382[17:29])
    OB Stepper_Y_M2_pad (.I(Stepper_Y_M2_c_2), .O(Stepper_Y_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(381[17:29])
    OB Stepper_Y_M1_pad (.I(Stepper_Y_M1_c_1), .O(Stepper_Y_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(380[17:29])
    OB Stepper_Y_M0_pad (.I(Stepper_Y_M0_c_0), .O(Stepper_Y_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(379[17:29])
    OB Stepper_Y_Dir_pad (.I(Stepper_Y_Dir_c), .O(Stepper_Y_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(378[17:30])
    OB Stepper_Y_Step_pad (.I(Stepper_Y_Step_c), .O(Stepper_Y_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(377[17:31])
    OB Stepper_X_En_pad (.I(Stepper_X_En_c), .O(Stepper_X_En));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(374[17:29])
    OB Stepper_X_M2_pad (.I(Stepper_X_M2_c_2), .O(Stepper_X_M2));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(373[17:29])
    OB Stepper_X_M1_pad (.I(Stepper_X_M1_c_1), .O(Stepper_X_M1));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(372[17:29])
    OB Stepper_X_M0_pad (.I(Stepper_X_M0_c_0), .O(Stepper_X_M0));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(371[17:29])
    OB Stepper_X_Dir_pad (.I(Stepper_X_Dir_c), .O(Stepper_X_Dir));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(370[17:30])
    OB Stepper_X_Step_pad (.I(Stepper_X_Step_c), .O(Stepper_X_Step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(369[17:31])
    OB status_led_pad_0 (.I(VCC_net), .O(status_led[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    OB status_led_pad_1 (.I(VCC_net), .O(status_led[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    LUT4 Select_3579_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[27]), 
         .D(n34317), .Z(n1)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3579_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3581_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[26]), 
         .D(n34317), .Z(n1_adj_398)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3581_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    OB status_led_pad_2 (.I(VCC_net), .O(status_led[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(366[20:30])
    OB uart_tx_pad (.I(n9395), .O(uart_tx));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(365[14:21])
    LUT4 Select_3583_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[25]), 
         .D(n34317), .Z(n1_adj_653)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3583_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3579_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[27]), 
         .D(rw), .Z(n2)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3579_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3585_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[24]), 
         .D(n34317), .Z(n1_adj_662)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3585_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3581_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[26]), 
         .D(rw), .Z(n2_adj_397)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3581_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3587_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[23]), 
         .D(n34317), .Z(n1_adj_666)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3587_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3589_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[22]), 
         .D(n34317), .Z(n1_adj_668)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3589_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3591_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[21]), 
         .D(n34317), .Z(n1_adj_646)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3591_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3593_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[20]), 
         .D(n34317), .Z(n1_adj_638)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3593_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_3_lut_rep_264_4_lut_4_lut (.A(n32439), .B(n30427), .C(n34317), 
         .D(prev_select_adj_559), .Z(n32358)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_rep_264_4_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n34320), .B(prev_select_adj_559), 
         .C(n30427), .D(n32439), .Z(n12620)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h1000;
    LUT4 i3_4_lut_rep_242 (.A(n54), .B(n6), .C(n1000), .D(n4_adj_598), 
         .Z(n32336)) /* synthesis lut_function=(!(A ((C)+!B)+!A ((C+!(D))+!B))) */ ;
    defparam i3_4_lut_rep_242.init = 16'h0c08;
    LUT4 Select_3583_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[25]), 
         .D(rw), .Z(n2_adj_651)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3583_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    FD1P3AX reset_count_2172_2173__i2 (.D(n66_adj_1129[1]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i2.GSR = "ENABLED";
    LUT4 LessThan_1434_i7_2_lut_rep_316 (.A(n7903[3]), .B(count_adj_845[3]), 
         .Z(n32410)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i7_2_lut_rep_316.init = 16'h6666;
    LUT4 i24631_4_lut (.A(n4), .B(n12), .C(n32352), .D(n30802), .Z(n14_adj_592)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24631_4_lut.init = 16'hcacc;
    LUT4 i8680_2_lut_3_lut (.A(n54), .B(n6), .C(n1000), .Z(n14446)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i8680_2_lut_3_lut.init = 16'h0808;
    LUT4 LessThan_1437_i4_4_lut (.A(count_adj_848[0]), .B(count_adj_848[1]), 
         .C(n7893[1]), .D(n7893[0]), .Z(n4)) /* synthesis lut_function=(A (B+!(C))+!A !(B (C (D))+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i4_4_lut.init = 16'h8ecf;
    LUT4 Select_3585_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[24]), 
         .D(rw), .Z(n2_adj_663)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3585_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3587_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[23]), 
         .D(rw), .Z(n2_adj_399)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3587_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i24629_4_lut (.A(n4_adj_616), .B(n12_adj_612), .C(n32356), .D(n30779), 
         .Z(n14_adj_611)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24629_4_lut.init = 16'hcacc;
    LUT4 Select_3589_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[22]), 
         .D(rw), .Z(n2_adj_667)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3589_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i24778_4_lut (.A(n32353), .B(n32352), .C(n32371), .D(n30797), 
         .Z(n30810)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24778_4_lut.init = 16'habaa;
    LUT4 i1_4_lut_adj_473 (.A(state_adj_834[5]), .B(state_adj_834[1]), .C(n183), 
         .D(n32), .Z(n15_adj_597)) /* synthesis lut_function=(!(A+!(B ((D)+!C)+!B !(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i1_4_lut_adj_473.init = 16'h4505;
    GSR GSR_INST (.GSR(VCC_net));
    FD1P3AX reset_count_2172_2173__i3 (.D(n66_adj_1129[2]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i3.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i4 (.D(n66_adj_1129[3]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i4.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i5 (.D(n66_adj_1129[4]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i5.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i6 (.D(n66_adj_1129[5]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i6.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i7 (.D(n66_adj_1129[6]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i7.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i8 (.D(n66_adj_1129[7]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i8.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i9 (.D(n66_adj_1129[8]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i9.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i10 (.D(n66_adj_1129[9]), .SP(n30), .CK(debug_c_c), 
            .Q(reset_count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i10.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i11 (.D(n66_adj_1129[10]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i11.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i12 (.D(n66_adj_1129[11]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i12.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i13 (.D(n66_adj_1129[12]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i13.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i14 (.D(n66_adj_1129[13]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i14.GSR = "ENABLED";
    FD1P3AX reset_count_2172_2173__i15 (.D(n66_adj_1129[14]), .SP(n30), 
            .CK(debug_c_c), .Q(reset_count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173__i15.GSR = "ENABLED";
    LUT4 i24637_2_lut (.A(bclk), .B(state_adj_834[1]), .Z(n30905)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(23[12:17])
    defparam i24637_2_lut.init = 16'h9999;
    LUT4 i24714_4_lut (.A(count_adj_845[9]), .B(count_adj_845[11]), .C(count_adj_845[12]), 
         .D(n6_adj_594), .Z(n28459)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i24714_4_lut.init = 16'h0001;
    LUT4 i24438_4_lut (.A(n32373), .B(n32399), .C(n32398), .D(n5_adj_648), 
         .Z(n30797)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24438_4_lut.init = 16'h5554;
    LUT4 LessThan_1434_i6_3_lut_3_lut (.A(n7903[3]), .B(count_adj_845[3]), 
         .C(count_adj_845[2]), .Z(n6_adj_614)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i6_3_lut_3_lut.init = 16'hd4d4;
    LUT4 Select_3591_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[21]), 
         .D(rw), .Z(n2_adj_593)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3591_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 LessThan_1437_i5_2_lut (.A(n7893[2]), .B(count_adj_848[2]), .Z(n5_adj_648)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i5_2_lut.init = 16'h6666;
    LUT4 i24665_4_lut (.A(n30457), .B(reset_count[14]), .C(n29618), .D(n19877), 
         .Z(n30)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam i24665_4_lut.init = 16'h373f;
    LUT4 i1_4_lut_adj_474 (.A(n20395), .B(n30456), .C(reset_count[6]), 
         .D(reset_count[5]), .Z(n30457)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[7:30])
    defparam i1_4_lut_adj_474.init = 16'hfcec;
    LUT4 i14656_4_lut (.A(reset_count[0]), .B(reset_count[4]), .C(n6_adj_396), 
         .D(reset_count[3]), .Z(n20395)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i14656_4_lut.init = 16'hccc8;
    LUT4 i2_2_lut (.A(reset_count[1]), .B(reset_count[2]), .Z(n6_adj_396)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1_2_lut (.A(reset_count[7]), .B(reset_count[8]), .Z(n30456)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(468[7:30])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(n32358), .B(n30423), .C(n34320), .Z(n12224)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i24722_4_lut_4_lut (.A(n32444), .B(n4_adj_519), .C(n9), .D(n1286[14]), 
         .Z(n12098)) /* synthesis lut_function=(!((B (C+!(D))+!B !(D))+!A)) */ ;
    defparam i24722_4_lut_4_lut.init = 16'h2a00;
    LUT4 i3_4_lut_4_lut (.A(n32444), .B(n32513), .C(n1286[8]), .D(n1286[0]), 
         .Z(n12788)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i3_4_lut_4_lut.init = 16'hfffd;
    LUT4 LessThan_1437_i7_2_lut_rep_304 (.A(n7893[3]), .B(count_adj_848[3]), 
         .Z(n32398)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i7_2_lut_rep_304.init = 16'h6666;
    LUT4 LessThan_1437_i6_3_lut_3_lut (.A(n7893[3]), .B(count_adj_848[3]), 
         .C(count_adj_848[2]), .Z(n6_adj_647)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i6_3_lut_3_lut.init = 16'hd4d4;
    LUT4 LessThan_1437_i9_2_lut_rep_305 (.A(n7893[4]), .B(count_adj_848[4]), 
         .Z(n32399)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i9_2_lut_rep_305.init = 16'h6666;
    LUT4 LessThan_1437_i8_3_lut_3_lut (.A(n7893[4]), .B(count_adj_848[4]), 
         .C(n6_adj_647), .Z(n8_adj_661)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1437_i8_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i2_3_lut_rep_260_4_lut_4_lut (.A(n34320), .B(n32443), .C(prev_select), 
         .D(n32401), .Z(n32354)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_rep_260_4_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_4_lut (.A(n34320), .B(register_addr[1]), .C(n32443), 
         .D(n32369), .Z(n30313)) /* synthesis lut_function=(A (B)+!A !((C (D))+!B)) */ ;
    defparam i1_2_lut_4_lut_4_lut.init = 16'h8ccc;
    LUT4 i13981_2_lut_2_lut (.A(n34320), .B(databus[4]), .Z(n580[4])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i13981_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_rep_256_3_lut_4_lut (.A(n32480), .B(n32439), .C(rw), 
         .D(prev_select), .Z(n32350)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_256_3_lut_4_lut.init = 16'h0004;
    LUT4 i24415_4_lut (.A(n32384), .B(n32411), .C(n32410), .D(n5_adj_615), 
         .Z(n30774)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam i24415_4_lut.init = 16'h5554;
    LUT4 LessThan_1434_i5_2_lut (.A(n7903[2]), .B(count_adj_845[2]), .Z(n5_adj_615)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i5_2_lut.init = 16'h6666;
    LUT4 Select_3621_i4_2_lut_3_lut_4_lut (.A(n32480), .B(n32439), .C(read_value_adj_695[4]), 
         .D(rw), .Z(n4_adj_617)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3621_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i24507_3_lut (.A(Stepper_A_M0_c_0), .B(stepping_adj_524), .C(register_addr[0]), 
         .Z(n30866)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24507_3_lut.init = 16'hcaca;
    LUT4 Select_3622_i4_2_lut_3_lut_4_lut (.A(n32480), .B(n32439), .C(read_value_adj_695[3]), 
         .D(n34317), .Z(n4_adj_607)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3622_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3623_i4_2_lut_3_lut_4_lut (.A(n32480), .B(n32439), .C(read_value_adj_695[2]), 
         .D(n34317), .Z(n4_adj_606)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3623_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i24508_3_lut (.A(div_factor_reg_adj_785[0]), .B(steps_reg_adj_786[0]), 
         .C(register_addr[0]), .Z(n30867)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24508_3_lut.init = 16'hcaca;
    LUT4 Select_3625_i4_2_lut_3_lut_4_lut (.A(n32480), .B(n32439), .C(read_value_adj_695[0]), 
         .D(rw), .Z(n4_adj_605)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3625_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3618_i4_2_lut_3_lut_4_lut (.A(n32480), .B(n32439), .C(read_value_adj_695[7]), 
         .D(rw), .Z(n4_adj_627)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3618_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3619_i4_2_lut_3_lut_4_lut (.A(n32480), .B(n32439), .C(read_value_adj_695[6]), 
         .D(rw), .Z(n4_adj_602)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3619_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3620_i4_2_lut_3_lut_4_lut (.A(n32480), .B(n32439), .C(read_value_adj_695[5]), 
         .D(rw), .Z(n4_adj_618)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3620_i4_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i13964_4_lut (.A(select[4]), .B(register_addr[5]), .C(n32454), 
         .D(register_addr[4]), .Z(arm_select[1])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(527[4] 556[11])
    defparam i13964_4_lut.init = 16'h0200;
    LUT4 Select_3593_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[20]), 
         .D(rw), .Z(n2_adj_639)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3593_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    VLO i1 (.Z(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i1_2_lut_rep_266_3_lut_4_lut (.A(n32505), .B(n32439), .C(rw), 
         .D(prev_select_adj_518), .Z(n32360)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_266_3_lut_4_lut.init = 16'h0004;
    LUT4 i2_3_lut_rep_272_4_lut_4_lut (.A(n34320), .B(n30240), .C(prev_select_adj_518), 
         .D(n32417), .Z(n32366)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_3_lut_rep_272_4_lut_4_lut.init = 16'h0100;
    LUT4 i14008_2_lut_2_lut (.A(n34320), .B(databus[0]), .Z(n571[0])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14008_2_lut_2_lut.init = 16'h4444;
    LUT4 LessThan_1434_i4_4_lut (.A(count_adj_845[0]), .B(count_adj_845[1]), 
         .C(n7903[1]), .D(n7903[0]), .Z(n4_adj_616)) /* synthesis lut_function=(A (B+!(C))+!A !(B (C (D))+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i4_4_lut.init = 16'h8ecf;
    LUT4 i14105_2_lut_2_lut (.A(n34320), .B(databus[2]), .Z(n580[2])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14105_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_4_lut_4_lut_adj_475 (.A(n34320), .B(register_addr[1]), 
         .C(n30240), .D(n32390), .Z(n30338)) /* synthesis lut_function=(A (B)+!A (B (C+!(D)))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_475.init = 16'hc8cc;
    GlobalControlPeripheral global_control (.n32448(n32448), .n32504(n32504), 
            .n11645(n11645), .register_addr({register_addr}), .read_value({read_value[31:2], 
            Open_0, read_value[0]}), .debug_c_c(debug_c_c), .n32379(n32379), 
            .n11753(n11753), .n30258(n30258), .n8048(n8048), .n21(n21_adj_600), 
            .n15(n15_adj_599), .read_size({read_size}), .n302(n302), .\register[2][0] (\register[2] [0]), 
            .n34321(n34321), .\register[0][2] (\register[0] [2]), .\select[1] (select[1]), 
            .n34323(n34323), .n34322(n34322), .\register[2][3] (\register[2] [3]), 
            .n28356(n28356), .n32422(n32422), .n32433(n32433), .n32429(n32429), 
            .n4(n4_adj_595), .n34317(n34317), .n32472(n32472), .rw(rw), 
            .n6(n6_adj_609), .force_pause(force_pause), .\databus[1] (databus[1]), 
            .n34320(n34320), .n20268(n20268), .xbee_pause_c(xbee_pause_c), 
            .n10513(n10513), .n14473(n14473), .signal_light_c(signal_light_c), 
            .\control_reg[7] (control_reg_adj_704[7]), .n28309(n28309), 
            .stepping(stepping), .n9633(n9633), .n14322(n14322), .\control_reg[7]_adj_188 (control_reg_adj_784[7]), 
            .n28270(n28270), .stepping_adj_189(stepping_adj_524), .\control_reg[7]_adj_190 (control_reg[7]), 
            .n28332(n28332), .n21_adj_191(n21), .\control_reg[7]_adj_192 (control_reg_adj_744[7]), 
            .n28296(n28296), .stepping_adj_193(stepping_adj_483), .n32503(n32503), 
            .n32455(n32455), .\select[4] (select[4]), .n32439(n32439), 
            .n32443(n32443), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(495[45] 505[74])
    \ArmPeripheral(axis_haddr=8'b0100000)  arm_z (.read_value({read_value_adj_747}), 
            .debug_c_c(debug_c_c), .n11981(n11981), .n32366(n32366), .\register_addr[1] (register_addr[1]), 
            .n30338(n30338), .\register_addr[0] (register_addr[0]), .Stepper_Z_M0_c_0(Stepper_Z_M0_c_0), 
            .stepping(stepping_adj_483), .VCC_net(VCC_net), .GND_net(GND_net), 
            .Stepper_Z_nFault_c(Stepper_Z_nFault_c), .n34322(n34322), .\read_size[0] (read_size_adj_748[0]), 
            .n30631(n30631), .n579(n571[0]), .prev_select(prev_select_adj_518), 
            .n32417(n32417), .n32505(n32505), .n32412(n32412), .n32390(n32390), 
            .rw(rw), .n34320(n34320), .n32360(n32360), .databus({databus}), 
            .n7852(n7852), .n34323(n34323), .n608(n580[4]), .n610(n580[2]), 
            .\control_reg[7] (control_reg_adj_744[7]), .Stepper_Z_En_c(Stepper_Z_En_c), 
            .n34324(n34324), .Stepper_Z_Dir_c(Stepper_Z_Dir_c), .Stepper_Z_M2_c_2(Stepper_Z_M2_c_2), 
            .Stepper_Z_M1_c_1(Stepper_Z_M1_c_1), .\read_size[2] (read_size_adj_748[2]), 
            .n29663(n29663), .\steps_reg[5] (steps_reg_adj_746[5]), .\steps_reg[3] (steps_reg_adj_746[3]), 
            .n34325(n34325), .n28296(n28296), .n14(n14_adj_650), .n15(n15_adj_669), 
            .n34317(n34317), .\register_addr[5] (register_addr[5]), .n30310(n30310), 
            .limit_c_2(limit_c_2), .\register_addr[4] (register_addr[4]), 
            .n32442(n32442), .n32503(n32503), .n32358(n32358), .n20505(n20505), 
            .Stepper_Z_Step_c(Stepper_Z_Step_c), .n32433(n32433)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(589[25] 602[45])
    \ArmPeripheral(axis_haddr=8'b0110000)  arm_a (.read_value({read_value_adj_787}), 
            .debug_c_c(debug_c_c), .n12620(n12620), .GND_net(GND_net), 
            .n30868(n30868), .register_addr({register_addr}), .n32504(n32504), 
            .n32503(n32503), .n30240(n30240), .\steps_reg[0] (steps_reg_adj_786[0]), 
            .n34323(n34323), .n3181({n3181}), .VCC_net(VCC_net), .Stepper_A_nFault_c(Stepper_A_nFault_c), 
            .\read_size[0] (read_size_adj_788[0]), .n30283(n30283), .Stepper_A_M0_c_0(Stepper_A_M0_c_0), 
            .n20505(n20505), .n579(n571[0]), .div_factor_reg({Open_1, 
            Open_2, Open_3, Open_4, Open_5, Open_6, Open_7, Open_8, 
            Open_9, Open_10, Open_11, Open_12, Open_13, Open_14, 
            Open_15, Open_16, Open_17, Open_18, Open_19, Open_20, 
            Open_21, Open_22, Open_23, Open_24, Open_25, Open_26, 
            Open_27, Open_28, Open_29, Open_30, Open_31, div_factor_reg_adj_785[0]}), 
            .n12224(n12224), .prev_select(prev_select_adj_559), .n32408(n32408), 
            .n32345(n32345), .n34321(n34321), .\databus[31] (databus[31]), 
            .\databus[28] (databus[28]), .n34322(n34322), .\databus[13] (databus[13]), 
            .\databus[11] (databus[11]), .\databus[10] (databus[10]), .\databus[9] (databus[9]), 
            .\databus[7] (databus[7]), .\databus[6] (databus[6]), .\databus[5] (databus[5]), 
            .n610(n580[2]), .\control_reg[7] (control_reg_adj_784[7]), .Stepper_A_En_c(Stepper_A_En_c), 
            .Stepper_A_Dir_c(Stepper_A_Dir_c), .\control_reg[4] (control_reg_adj_784[4]), 
            .\databus[4] (databus[4]), .\databus[3] (databus[3]), .Stepper_A_M2_c_2(Stepper_A_M2_c_2), 
            .Stepper_A_M1_c_1(Stepper_A_M1_c_1), .\databus[1] (databus[1]), 
            .\read_size[2] (read_size_adj_788[2]), .n30284(n30284), .n34324(n34324), 
            .n34325(n34325), .\steps_reg[16] (steps_reg_adj_786[16]), .\steps_reg[8] (steps_reg_adj_786[8]), 
            .\steps_reg[5] (steps_reg_adj_786[5]), .\steps_reg[4] (steps_reg_adj_786[4]), 
            .\steps_reg[3] (steps_reg_adj_786[3]), .n32360(n32360), .n7852(n7852), 
            .\register[0][2] (\register[0] [2]), .force_pause(force_pause), 
            .n21(n21_adj_600), .n32480(n32480), .n32481(n32481), .n32440(n32440), 
            .n32412(n32412), .n6124(n6096[4]), .n30211(n30211), .n17(n17), 
            .n224({n224_adj_791}), .stepping(stepping_adj_524), .n34320(n34320), 
            .n32454(n32454), .\register[2][0] (\register[2] [0]), .n15(n15_adj_599), 
            .\register[2][3] (\register[2] [3]), .n4(n4_adj_595), .n32460(n32460), 
            .n32442(n32442), .\div_factor_reg[4] (div_factor_reg_adj_785[4]), 
            .\div_factor_reg[8] (div_factor_reg_adj_785[8]), .\databus[8] (databus[8]), 
            .\databus[12] (databus[12]), .\databus[14] (databus[14]), .\databus[15] (databus[15]), 
            .\div_factor_reg[16] (div_factor_reg_adj_785[16]), .\databus[16] (databus[16]), 
            .\databus[17] (databus[17]), .\databus[18] (databus[18]), .\databus[19] (databus[19]), 
            .\databus[20] (databus[20]), .\databus[21] (databus[21]), .\databus[22] (databus[22]), 
            .\databus[23] (databus[23]), .\databus[24] (databus[24]), .\databus[25] (databus[25]), 
            .\databus[26] (databus[26]), .\databus[27] (databus[27]), .\databus[29] (databus[29]), 
            .\databus[30] (databus[30]), .limit_c_3(limit_c_3), .Stepper_A_Step_c(Stepper_A_Step_c), 
            .n15_adj_187(n15_adj_395), .n28270(n28270), .n14(n14), .n32381(n32381), 
            .n30427(n30427), .rw(rw), .n32433(n32433)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(604[25] 617[45])
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_476 (.A(n34320), .B(prev_select_adj_518), 
         .C(n32439), .D(n32505), .Z(n11981)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_476.init = 16'h0010;
    LUT4 Select_3624_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[1]), 
         .D(rw), .Z(n1_adj_608)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3624_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 LessThan_1434_i13_2_lut_rep_289 (.A(n7903[6]), .B(count_adj_845[6]), 
         .Z(n32383)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i13_2_lut_rep_289.init = 16'h6666;
    \ArmPeripheral(axis_haddr=8'b010000)  arm_y (.databus({databus}), .n3363(n3363), 
            .debug_c_c(debug_c_c), .n34322(n34322), .VCC_net(VCC_net), 
            .GND_net(GND_net), .Stepper_Y_nFault_c(Stepper_Y_nFault_c), 
            .\read_size[0] (read_size_adj_708[0]), .n30710(n30710), .Stepper_Y_M0_c_0(Stepper_Y_M0_c_0), 
            .n579(n571[0]), .\register_addr[5] (register_addr[5]), .\register_addr[4] (register_addr[4]), 
            .n11883(n11883), .n12434(n12434), .\arm_select[1] (arm_select[1]), 
            .read_value({read_value_adj_707}), .n32504(n32504), .n32503(n32503), 
            .n32480(n32480), .\select[4] (select[4]), .n32401(n32401), 
            .n32348(n32348), .n34321(n34321), .n34324(n34324), .n34323(n34323), 
            .n34325(n34325), .\control_reg[7] (control_reg_adj_704[7]), 
            .Stepper_Y_En_c(Stepper_Y_En_c), .Stepper_Y_Dir_c(Stepper_Y_Dir_c), 
            .Stepper_Y_M2_c_2(Stepper_Y_M2_c_2), .Stepper_Y_M1_c_1(Stepper_Y_M1_c_1), 
            .\read_size[2] (read_size_adj_708[2]), .n30411(n30411), .n30427(n30427), 
            .n32408(n32408), .n32505(n32505), .n32417(n32417), .n34326(n34326), 
            .\steps_reg[5] (steps_reg_adj_706[5]), .\steps_reg[3] (steps_reg_adj_706[3]), 
            .limit_c_1(limit_c_1), .stepping(stepping), .\register_addr[0] (register_addr[0]), 
            .n34320(n34320), .\register_addr[1] (register_addr[1]), .n14(n14_adj_665), 
            .n15(n15_adj_400), .n28309(n28309), .n32412(n32412), .n32389(n32389), 
            .rw(rw), .Stepper_Y_Step_c(Stepper_Y_Step_c), .n52(n52), .n34317(n34317), 
            .n32365(n32365), .n32433(n32433)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(574[25] 587[45])
    LUT4 Select_3601_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[16]), 
         .D(rw), .Z(n1_adj_644)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3601_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3595_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[19]), 
         .D(rw), .Z(n2_adj_635)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3595_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3599_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[17]), 
         .D(rw), .Z(n2_adj_637)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3599_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_477 (.A(n34320), .B(prev_select), 
         .C(n32439), .D(n32480), .Z(n11966)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_477.init = 16'h0010;
    RCPeripheral rc_receiver (.\read_value[13] (read_value[13]), .n1(n1_adj_630), 
            .n32472(n32472), .\read_value[13]_adj_43 (read_value_adj_695[13]), 
            .read_value({read_value_adj_707}), .n32375(n32375), .n52(n52), 
            .\register_addr[0] (register_addr[0]), .databus_out({databus_out}), 
            .n2(n2_adj_629), .rw(rw), .databus({databus}), .\read_value[12]_adj_45 (read_value[12]), 
            .n1_adj_46(n1_adj_628), .n4(n4_adj_606), .\read_value[12]_adj_47 (read_value_adj_695[12]), 
            .n2_adj_48(n2_adj_624), .\read_value[11]_adj_49 (read_value[11]), 
            .n1_adj_50(n1_adj_623), .\read_value[11]_adj_51 (read_value_adj_695[11]), 
            .\select[7] (select[7]), .n32504(n32504), .n32481(n32481), 
            .\register_addr[1] (register_addr[1]), .n30427(n30427), .n30283(n30283), 
            .n30284(n30284), .n32505(n32505), .n30631(n30631), .n29663(n29663), 
            .n11883(n11883), .n30710(n30710), .n30411(n30411), .n2_adj_52(n2_adj_620), 
            .\read_value[10]_adj_53 (read_value[10]), .n1_adj_54(n1_adj_619), 
            .\read_value[10]_adj_55 (read_value_adj_695[10]), .\register_addr[4] (register_addr[4]), 
            .\read_size[0] (read_size_adj_696[0]), .\read_size[0]_adj_56 (read_size_adj_748[0]), 
            .\register_addr[5] (register_addr[5]), .\read_size[0]_adj_57 (read_size_adj_708[0]), 
            .\read_size[0]_adj_58 (read_size_adj_788[0]), .n2_adj_59(n2_adj_641), 
            .n2_adj_60(n2_adj_663), .\read_value[18]_adj_61 (read_value[18]), 
            .n1_adj_62(n1_adj_640), .\read_value[18]_adj_63 (read_value_adj_695[18]), 
            .\read_value[2]_adj_64 (read_value_adj_787[2]), .n32374(n32374), 
            .\read_value[24]_adj_65 (read_value[24]), .n1_adj_66(n1_adj_662), 
            .n2_adj_67(n2_adj_626), .\read_value[2]_adj_68 (read_value_adj_747[2]), 
            .\read_value[2]_adj_69 (read_value[2]), .n32376(n32376), .\read_value[9]_adj_70 (read_value[9]), 
            .n1_adj_71(n1_adj_625), .\read_value[24]_adj_72 (read_value_adj_695[24]), 
            .\read_value[9]_adj_73 (read_value_adj_695[9]), .n32455(n32455), 
            .\register_addr[2] (register_addr[2]), .\register_addr[3] (register_addr[3]), 
            .n30401(n30401), .read_value_adj_186({read_value_adj_690}), 
            .n64(n64), .n2_adj_82(n2_adj_637), .\read_value[17]_adj_83 (read_value[17]), 
            .n1_adj_84(n1_adj_636), .\read_value[17]_adj_85 (read_value_adj_695[17]), 
            .n2_adj_86(n2_adj_399), .n2_adj_87(n2_adj_645), .\read_value[16]_adj_88 (read_value[16]), 
            .n1_adj_89(n1_adj_644), .\read_value[16]_adj_90 (read_value_adj_695[16]), 
            .read_size({read_size}), .\select[1] (select[1]), .n32486(n32486), 
            .\sendcount[1] (sendcount[1]), .n11271(n11271), .n2_adj_92(n2_adj_643), 
            .\read_value[15]_adj_93 (read_value[15]), .n1_adj_94(n1_adj_642), 
            .n2_adj_95(n2_adj_622), .\read_value[15]_adj_96 (read_value_adj_695[15]), 
            .\read_value[23]_adj_97 (read_value[23]), .n1_adj_98(n1_adj_666), 
            .n32381(n32381), .n30423(n30423), .n32345(n32345), .\read_value[8]_adj_99 (read_value[8]), 
            .n1_adj_100(n1_adj_621), .n1_adj_101(n1_adj_608), .n2_adj_102(n2_adj_633), 
            .\read_value[14]_adj_103 (read_value[14]), .n1_adj_104(n1_adj_632), 
            .\read_value[8]_adj_105 (read_value_adj_695[8]), .\read_value[14]_adj_106 (read_value_adj_695[14]), 
            .\read_value[1]_adj_107 (read_value_adj_695[1]), .n6(n6_adj_609), 
            .\read_value[23]_adj_108 (read_value_adj_695[23]), .n2_adj_109(n2_adj_631), 
            .\read_value[1]_adj_110 (read_value_adj_747[1]), .n2_adj_111(n2_adj_667), 
            .\read_value[22]_adj_112 (read_value[22]), .n1_adj_113(n1_adj_668), 
            .\read_value[22]_adj_114 (read_value_adj_695[22]), .n2_adj_115(n2_adj_601), 
            .n2_adj_116(n2_adj_635), .\read_value[30]_adj_117 (read_value[30]), 
            .n1_adj_118(n1_adj_649), .\read_value[19]_adj_119 (read_value[19]), 
            .n1_adj_120(n1_adj_634), .n4_adj_121(n4_adj_627), .\read_value[7]_adj_122 (read_value_adj_787[7]), 
            .\read_value[30]_adj_123 (read_value_adj_695[30]), .n2_adj_124(n2_adj_664), 
            .\read_value[19]_adj_125 (read_value_adj_695[19]), .\read_size[2]_adj_126 (read_size_adj_696[2]), 
            .\read_size[2]_adj_127 (read_size_adj_748[2]), .\read_size[2]_adj_128 (read_size_adj_708[2]), 
            .\read_size[2]_adj_129 (read_size_adj_788[2]), .\read_value[7]_adj_130 (read_value_adj_747[7]), 
            .\read_value[7]_adj_131 (read_value[7]), .n34317(n34317), .\read_value[29]_adj_132 (read_value[29]), 
            .n1_adj_133(n1_adj_520), .n2_adj_134(n2_adj_593), .n4_adj_135(n4_adj_602), 
            .\read_value[6]_adj_136 (read_value_adj_787[6]), .\read_value[6]_adj_137 (read_value_adj_747[6]), 
            .\read_value[6]_adj_138 (read_value[6]), .\read_value[29]_adj_139 (read_value_adj_695[29]), 
            .n4_adj_140(n4_adj_605), .\read_value[0]_adj_141 (read_value_adj_787[0]), 
            .\read_value[0]_adj_142 (read_value_adj_747[0]), .\read_value[0]_adj_143 (read_value[0]), 
            .\read_value[21]_adj_144 (read_value[21]), .n1_adj_145(n1_adj_646), 
            .n4_adj_146(n4_adj_618), .\read_value[5]_adj_147 (read_value_adj_787[5]), 
            .\read_value[5]_adj_148 (read_value_adj_747[5]), .\read_value[5]_adj_149 (read_value[5]), 
            .\read_value[21]_adj_150 (read_value_adj_695[21]), .n2_adj_151(n2_adj_639), 
            .\select[2] (select[2]), .\read_size[0]_adj_152 (read_size_adj_691[0]), 
            .n5(n5), .n32439(n32439), .n6_adj_153(n6_adj_596), .n2_adj_154(n2_adj_603), 
            .\read_value[31]_adj_155 (read_value[31]), .n1_adj_156(n1_adj_604), 
            .\read_value[31]_adj_157 (read_value_adj_695[31]), .\reg_size[2] (reg_size[2]), 
            .n2_adj_158(n2_adj_444), .\read_value[28]_adj_159 (read_value[28]), 
            .n1_adj_160(n1_adj_652), .\read_value[28]_adj_161 (read_value_adj_695[28]), 
            .\read_value[20]_adj_162 (read_value[20]), .n1_adj_163(n1_adj_638), 
            .n4_adj_164(n4_adj_617), .\read_value[4]_adj_165 (read_value_adj_787[4]), 
            .\read_value[4]_adj_166 (read_value_adj_747[4]), .\read_value[4]_adj_167 (read_value[4]), 
            .\read_value[20]_adj_168 (read_value_adj_695[20]), .n2_adj_169(n2), 
            .\read_value[27]_adj_170 (read_value[27]), .n1_adj_171(n1), 
            .\read_value[27]_adj_172 (read_value_adj_695[27]), .n2_adj_173(n2_adj_397), 
            .\read_value[26]_adj_174 (read_value[26]), .n1_adj_175(n1_adj_398), 
            .\read_value[26]_adj_176 (read_value_adj_695[26]), .n4_adj_177(n4_adj_607), 
            .\read_value[3]_adj_178 (read_value_adj_787[3]), .\read_value[3]_adj_179 (read_value_adj_747[3]), 
            .\read_value[3]_adj_180 (read_value[3]), .n2_adj_181(n2_adj_651), 
            .\read_value[25]_adj_182 (read_value[25]), .n1_adj_183(n1_adj_653), 
            .\read_value[25]_adj_184 (read_value_adj_695[25]), .debug_c_c(debug_c_c), 
            .n28324(n28324), .GND_net(GND_net), .n32341(n32341), .rc_ch8_c(rc_ch8_c), 
            .n31024(n31024), .n30913(n30913), .n12030(n12030), .n31005(n31005), 
            .n28308(n28308), .rc_ch7_c(rc_ch7_c), .n30995(n30995), .n12031(n12031), 
            .n30929(n30929), .rc_ch4_c(rc_ch4_c), .n28304(n28304), .n12138(n12138), 
            .n31000(n31000), .n30969(n30969), .n28317(n28317), .rc_ch3_c(rc_ch3_c), 
            .n1000(n1000), .n988(n988), .n32336(n32336), .n14446(n14446), 
            .rc_ch2_c(rc_ch2_c), .n54(n54), .n4_adj_185(n4_adj_598), .n12841(n12841), 
            .n31049(n31049), .n28312(n28312), .rc_ch1_c(rc_ch1_c), .n30911(n30911)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(622[15] 634[41])
    LUT4 Select_3599_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[17]), 
         .D(rw), .Z(n1_adj_636)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3599_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 Select_3601_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[16]), 
         .D(rw), .Z(n2_adj_645)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3601_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 Select_3597_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[18]), 
         .D(rw), .Z(n2_adj_641)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3597_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 LessThan_1434_i10_3_lut_3_lut (.A(n7903[6]), .B(count_adj_845[6]), 
         .C(count_adj_845[5]), .Z(n10_adj_613)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[9:43])
    defparam LessThan_1434_i10_3_lut_3_lut.init = 16'hd4d4;
    \ProtocolInterface(baud_div=12)  protocol_interface (.debug_c_c(debug_c_c), 
            .register_addr({register_addr}), .n32389(n32389), .n30258(n30258), 
            .n3363(n3363), .n30423(n30423), .n32348(n32348), .n1318(n1286[0]), 
            .n1304(n1286[14]), .n1310(n1286[8]), .n12098(n12098), .databus_out({databus_out}), 
            .n32444(n32444), .n32358(n32358), .databus({databus}), .n224({n224_adj_791}), 
            .n3181({n3181}), .\select[1] (select[1]), .n12788(n12788), 
            .\sendcount[1] (sendcount[1]), .debug_c_7(debug_c_7), .\select[2] (select[2]), 
            .\select[4] (select[4]), .\select[7] (select[7]), .\steps_reg[4] (steps_reg_adj_786[4]), 
            .n15(n15), .n9(n9), .n30310(n30310), .n32343(n32343), .n224_adj_42({n224}), 
            .n3451({n3451}), .\steps_reg[7] (steps_reg[7]), .n13(n13), 
            .\steps_reg[3] (steps_reg_adj_786[3]), .n15_adj_33(n15_adj_395), 
            .rw(rw), .\steps_reg[5] (steps_reg_adj_786[5]), .n14(n14), 
            .n4(n4_adj_519), .n34317(n34317), .\steps_reg[5]_adj_34 (steps_reg_adj_706[5]), 
            .n14_adj_35(n14_adj_665), .\steps_reg[3]_adj_36 (steps_reg_adj_706[3]), 
            .n15_adj_37(n15_adj_400), .\steps_reg[5]_adj_38 (steps_reg_adj_746[5]), 
            .n14_adj_39(n14_adj_650), .\steps_reg[3]_adj_40 (steps_reg_adj_746[3]), 
            .n15_adj_41(n15_adj_669), .n32513(n32513), .n11271(n11271), 
            .n5(n5), .n6(n6_adj_596), .\reg_size[2] (reg_size[2]), .n32486(n32486), 
            .debug_c_2(debug_c_2), .debug_c_3(debug_c_3), .debug_c_4(debug_c_4), 
            .debug_c_5(debug_c_5), .n34320(n34320), .n32503(n32503), .n30401(n30401), 
            .n11753(n11753), .\reset_count[14] (reset_count[14]), .\reset_count[12] (reset_count[12]), 
            .\reset_count[13] (reset_count[13]), .\reset_count[11] (reset_count[11]), 
            .n19877(n19877), .\reset_count[8] (reset_count[8]), .n27962(n27962), 
            .n9395(n9395), .\reset_count[10] (reset_count[10]), .\reset_count[9] (reset_count[9]), 
            .GND_net(GND_net), .state({state_adj_834}), .n32(n32), .\rdata[0] (rdata[0]), 
            .bclk(bclk), .n29158(n29158), .\rdata[1] (rdata[1]), .n9396_c(n9396_c), 
            .n31442(n31442), .n183(n183), .n31427(n31427), .n32432(n32432), 
            .n32409(n32409), .n32495(n32495), .n32494(n32494)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(475[26] 485[57])
    LUT4 Select_3603_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[15]), 
         .D(rw), .Z(n2_adj_643)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3603_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    \ArmPeripheral(axis_haddr=8'b0)  arm_x (.\register_addr[0] (register_addr[0]), 
            .debug_c_c(debug_c_c), .n34324(n34324), .n3451({n3451}), .n32401(n32401), 
            .prev_select(prev_select), .\register_addr[5] (register_addr[5]), 
            .n34317(n34317), .n32343(n32343), .n34321(n34321), .limit_c_0(limit_c_0), 
            .n32481(n32481), .n32480(n32480), .n32460(n32460), .n302(n302), 
            .\register_addr[1] (register_addr[1]), .n32504(n32504), .n30726(n30726), 
            .n32422(n32422), .\read_size[0] (read_size_adj_696[0]), .n11966(n11966), 
            .n34322(n34322), .Stepper_X_M0_c_0(Stepper_X_M0_c_0), .n579(n571[0]), 
            .n34323(n34323), .\steps_reg[7] (steps_reg[7]), .read_value({read_value_adj_695}), 
            .\databus[31] (databus[31]), .n34325(n34325), .\databus[30] (databus[30]), 
            .\databus[29] (databus[29]), .\databus[26] (databus[26]), .\databus[13] (databus[13]), 
            .\databus[11] (databus[11]), .\databus[10] (databus[10]), .\databus[9] (databus[9]), 
            .\databus[7] (databus[7]), .\databus[6] (databus[6]), .\databus[5] (databus[5]), 
            .n608(n580[4]), .n610(n580[2]), .\control_reg[7] (control_reg[7]), 
            .Stepper_X_En_c(Stepper_X_En_c), .n34326(n34326), .Stepper_X_Dir_c(Stepper_X_Dir_c), 
            .\databus[3] (databus[3]), .Stepper_X_M2_c_2(Stepper_X_M2_c_2), 
            .Stepper_X_M1_c_1(Stepper_X_M1_c_1), .\databus[1] (databus[1]), 
            .\read_size[2] (read_size_adj_696[2]), .n32433(n32433), .\register_addr[4] (register_addr[4]), 
            .\register_addr[3] (register_addr[3]), .n11753(n11753), .n30310(n30310), 
            .n30313(n30313), .n11645(n11645), .n34320(n34320), .GND_net(GND_net), 
            .n224({n224}), .n21(n21), .n30423(n30423), .n32365(n32365), 
            .n12434(n12434), .\register_addr[6] (register_addr[6]), .\register_addr[7] (register_addr[7]), 
            .n32448(n32448), .n32503(n32503), .n20268(n20268), .n28356(n28356), 
            .\databus[8] (databus[8]), .\databus[12] (databus[12]), .\databus[14] (databus[14]), 
            .\databus[15] (databus[15]), .n32455(n32455), .n32442(n32442), 
            .n32369(n32369), .rw(rw), .n32350(n32350), .\databus[16] (databus[16]), 
            .\databus[17] (databus[17]), .\databus[18] (databus[18]), .\databus[19] (databus[19]), 
            .\databus[20] (databus[20]), .\databus[21] (databus[21]), .\databus[22] (databus[22]), 
            .\databus[23] (databus[23]), .n32354(n32354), .\databus[24] (databus[24]), 
            .\databus[25] (databus[25]), .\databus[27] (databus[27]), .\databus[28] (databus[28]), 
            .VCC_net(VCC_net), .Stepper_X_nFault_c(Stepper_X_nFault_c), 
            .n28332(n28332), .n32379(n32379), .n30401(n30401), .n8048(n8048), 
            .n13(n13), .Stepper_X_Step_c(Stepper_X_Step_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(559[25] 572[45])
    CCU2D reset_count_2172_2173_add_4_15 (.A0(reset_count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27764), .S0(n66_adj_1129[13]), 
          .S1(n66_adj_1129[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_15.INIT0 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_15.INIT1 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_15.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_15.INJECT1_1 = "NO";
    CCU2D reset_count_2172_2173_add_4_13 (.A0(reset_count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27763), .COUT(n27764), .S0(n66_adj_1129[11]), 
          .S1(n66_adj_1129[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_13.INIT0 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_13.INIT1 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_13.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_13.INJECT1_1 = "NO";
    CCU2D reset_count_2172_2173_add_4_11 (.A0(reset_count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27762), .COUT(n27763), .S0(n66_adj_1129[9]), 
          .S1(n66_adj_1129[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_11.INIT0 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_11.INIT1 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_11.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_11.INJECT1_1 = "NO";
    CCU2D reset_count_2172_2173_add_4_9 (.A0(reset_count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27761), .COUT(n27762), .S0(n66_adj_1129[7]), 
          .S1(n66_adj_1129[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_9.INIT0 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_9.INIT1 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_9.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_9.INJECT1_1 = "NO";
    CCU2D reset_count_2172_2173_add_4_7 (.A0(reset_count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27760), .COUT(n27761), .S0(n66_adj_1129[5]), 
          .S1(n66_adj_1129[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_7.INIT0 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_7.INIT1 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_7.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_7.INJECT1_1 = "NO";
    LUT4 Select_3605_i2_2_lut_3_lut_4_lut (.A(n32505), .B(n32439), .C(read_value_adj_747[14]), 
         .D(rw), .Z(n2_adj_633)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam Select_3605_i2_2_lut_3_lut_4_lut.init = 16'h4000;
    CCU2D reset_count_2172_2173_add_4_5 (.A0(reset_count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27759), .COUT(n27760), .S0(n66_adj_1129[3]), 
          .S1(n66_adj_1129[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_5.INIT0 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_5.INIT1 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_5.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_5.INJECT1_1 = "NO";
    CCU2D reset_count_2172_2173_add_4_3 (.A0(reset_count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(reset_count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27758), .COUT(n27759), .S0(n66_adj_1129[1]), 
          .S1(n66_adj_1129[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_3.INIT0 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_3.INIT1 = 16'hfaaa;
    defparam reset_count_2172_2173_add_4_3.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_3.INJECT1_1 = "NO";
    CCU2D reset_count_2172_2173_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(reset_count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27758), .S1(n66_adj_1129[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(469[20:35])
    defparam reset_count_2172_2173_add_4_1.INIT0 = 16'hF000;
    defparam reset_count_2172_2173_add_4_1.INIT1 = 16'h0555;
    defparam reset_count_2172_2173_add_4_1.INJECT1_0 = "NO";
    defparam reset_count_2172_2173_add_4_1.INJECT1_1 = "NO";
    ClockDivider_U10 pwm_clk_div (.debug_c_c(debug_c_c), .n241(n241), .n34320(n34320), 
            .n6674(n6674), .n32341(n32341), .n30913(n30913), .n12030(n12030), 
            .n30995(n30995), .n12031(n12031), .n30929(n30929), .n28304(n28304), 
            .n30911(n30911), .n28312(n28312), .n31000(n31000), .n28317(n28317), 
            .n31005(n31005), .n28308(n28308), .n31024(n31024), .n28324(n28324), 
            .n988(n988), .n6(n6), .n31049(n31049), .n12841(n12841), 
            .n30969(n30969), .n12138(n12138), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(508[15] 511[41])
    LUT4 Select_3597_i1_2_lut_3_lut_4_lut (.A(n32439), .B(n30427), .C(read_value_adj_787[18]), 
         .D(rw), .Z(n1_adj_640)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam Select_3597_i1_2_lut_3_lut_4_lut.init = 16'h8000;
    
endmodule
//
// Verilog Description of module PWMPeripheral
//

module PWMPeripheral (\read_size[0] , debug_c_c, n30726, n34322, \databus[0] , 
            \select[2] , rw, n32440, \register_addr[0] , read_value, 
            n282, n34326, \databus[6] , \databus[5] , \databus[4] , 
            \databus[3] , \databus[2] , \databus[1] , n32448, n32460, 
            n34320, n34317, n64, \count[0] , n32341, motor_pwm_r_c, 
            GND_net, n9633, n14322, \count[1] , \count[2] , \count[3] , 
            \count[4] , \count[5] , \count[6] , \count[7] , \count[8] , 
            n3589, n7893, n7902, n10513, n14473, \count[0]_adj_195 , 
            \count[12] , \count[11] , \count[9] , \count[8]_adj_196 , 
            \count[6]_adj_197 , \count[5]_adj_198 , \count[3]_adj_199 , 
            \count[2]_adj_200 , \count[1]_adj_201 , motor_pwm_l_c, n28459, 
            n32356, n10, n12, \reset_count[6] , n30456, \reset_count[4] , 
            \reset_count[5] , n30458, \reset_count[12] , \reset_count[11] , 
            \reset_count[13] , n29618, n3586, n6, n32411, n6_adj_202, 
            n8, n7912, n7906, n7905, n7908, n7910, n7909, n7911) /* synthesis syn_module_defined=1 */ ;
    output \read_size[0] ;
    input debug_c_c;
    input n30726;
    input n34322;
    input \databus[0] ;
    input \select[2] ;
    input rw;
    input n32440;
    input \register_addr[0] ;
    output [7:0]read_value;
    input n282;
    input n34326;
    input \databus[6] ;
    input \databus[5] ;
    input \databus[4] ;
    input \databus[3] ;
    input \databus[2] ;
    input \databus[1] ;
    input n32448;
    input n32460;
    input n34320;
    input n34317;
    output n64;
    output \count[0] ;
    input n32341;
    output motor_pwm_r_c;
    input GND_net;
    output n9633;
    input n14322;
    output \count[1] ;
    output \count[2] ;
    output \count[3] ;
    output \count[4] ;
    output \count[5] ;
    output \count[6] ;
    output \count[7] ;
    output \count[8] ;
    input n3589;
    output [7:0]n7893;
    output n7902;
    output n10513;
    input n14473;
    output \count[0]_adj_195 ;
    output \count[12] ;
    output \count[11] ;
    output \count[9] ;
    output \count[8]_adj_196 ;
    output \count[6]_adj_197 ;
    output \count[5]_adj_198 ;
    output \count[3]_adj_199 ;
    output \count[2]_adj_200 ;
    output \count[1]_adj_201 ;
    output motor_pwm_l_c;
    input n28459;
    output n32356;
    input n10;
    output n12;
    input \reset_count[6] ;
    input n30456;
    input \reset_count[4] ;
    input \reset_count[5] ;
    output n30458;
    input \reset_count[12] ;
    input \reset_count[11] ;
    input \reset_count[13] ;
    output n29618;
    input n3586;
    output n6;
    output n32411;
    input n6_adj_202;
    output n8;
    output n7912;
    output n7906;
    output n7905;
    output n7908;
    output n7910;
    output n7909;
    output n7911;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n12099;
    wire [7:0]\register[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(55[12:20])
    
    wire n32392, prev_select, n32511, n32394, n8052;
    wire [7:0]n4894;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(55[12:20])
    
    wire n12566, n20489, n32418;
    
    FD1P3AX read_size__i1 (.D(n30726), .SP(n12099), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3JX register_0__i1 (.D(\databus[0] ), .SP(n32392), .PD(n34322), 
            .CK(debug_c_c), .Q(\register[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i1.GSR = "ENABLED";
    FD1S3AX prev_select_138 (.D(\select[2] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam prev_select_138.GSR = "ENABLED";
    LUT4 i3870_2_lut_rep_300_4_lut (.A(rw), .B(n32511), .C(n32440), .D(\register_addr[0] ), 
         .Z(n32394)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i3870_2_lut_rep_300_4_lut.init = 16'h0400;
    FD1P3IX read_value__i1 (.D(n4894[1]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n4894[2]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n4894[3]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n4894[4]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n4894[5]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3AX register_0__i16 (.D(n282), .SP(n12566), .CK(debug_c_c), .Q(\register[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i16.GSR = "ENABLED";
    FD1P3JX register_0__i15 (.D(\databus[6] ), .SP(n32394), .PD(n34326), 
            .CK(debug_c_c), .Q(\register[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i15.GSR = "ENABLED";
    FD1P3JX register_0__i14 (.D(\databus[5] ), .SP(n32394), .PD(n34326), 
            .CK(debug_c_c), .Q(\register[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i14.GSR = "ENABLED";
    FD1P3JX register_0__i13 (.D(\databus[4] ), .SP(n32394), .PD(n34326), 
            .CK(debug_c_c), .Q(\register[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i13.GSR = "ENABLED";
    FD1P3JX register_0__i12 (.D(\databus[3] ), .SP(n32394), .PD(n34326), 
            .CK(debug_c_c), .Q(\register[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i12.GSR = "ENABLED";
    FD1P3JX register_0__i11 (.D(\databus[2] ), .SP(n32394), .PD(n34326), 
            .CK(debug_c_c), .Q(\register[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i11.GSR = "ENABLED";
    FD1P3JX register_0__i10 (.D(\databus[1] ), .SP(n32394), .PD(n34326), 
            .CK(debug_c_c), .Q(\register[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i10.GSR = "ENABLED";
    FD1P3JX register_0__i9 (.D(\databus[0] ), .SP(n32394), .PD(n34326), 
            .CK(debug_c_c), .Q(\register[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i9.GSR = "ENABLED";
    FD1P3AX register_0__i8 (.D(n282), .SP(n20489), .CK(debug_c_c), .Q(\register[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i8.GSR = "ENABLED";
    FD1P3JX register_0__i7 (.D(\databus[6] ), .SP(n32392), .PD(n34326), 
            .CK(debug_c_c), .Q(\register[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i7.GSR = "ENABLED";
    FD1P3JX register_0__i6 (.D(\databus[5] ), .SP(n32392), .PD(n34326), 
            .CK(debug_c_c), .Q(\register[0] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i6.GSR = "ENABLED";
    FD1P3JX register_0__i5 (.D(\databus[4] ), .SP(n32392), .PD(n34326), 
            .CK(debug_c_c), .Q(\register[0] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i5.GSR = "ENABLED";
    FD1P3JX register_0__i4 (.D(\databus[3] ), .SP(n32392), .PD(n34326), 
            .CK(debug_c_c), .Q(\register[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i4.GSR = "ENABLED";
    FD1P3JX register_0__i3 (.D(\databus[2] ), .SP(n32392), .PD(n34326), 
            .CK(debug_c_c), .Q(\register[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i3.GSR = "ENABLED";
    FD1P3JX register_0__i2 (.D(\databus[1] ), .SP(n32392), .PD(n34326), 
            .CK(debug_c_c), .Q(\register[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam register_0__i2.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n4894[6]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n4894[7]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i7.GSR = "ENABLED";
    LUT4 mux_1586_Mux_1_i1_3_lut (.A(\register[0] [1]), .B(\register[1] [1]), 
         .C(\register_addr[0] ), .Z(n4894[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1586_Mux_2_i1_3_lut (.A(\register[0] [2]), .B(\register[1] [2]), 
         .C(\register_addr[0] ), .Z(n4894[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1586_Mux_3_i1_3_lut (.A(\register[0] [3]), .B(\register[1] [3]), 
         .C(\register_addr[0] ), .Z(n4894[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1586_Mux_4_i1_3_lut (.A(\register[0] [4]), .B(\register[1] [4]), 
         .C(\register_addr[0] ), .Z(n4894[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_4_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1586_Mux_5_i1_3_lut (.A(\register[0] [5]), .B(\register[1] [5]), 
         .C(\register_addr[0] ), .Z(n4894[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_5_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1586_Mux_6_i1_3_lut (.A(\register[0] [6]), .B(\register[1] [6]), 
         .C(\register_addr[0] ), .Z(n4894[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_6_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1586_Mux_7_i1_3_lut (.A(\register[0] [7]), .B(\register[1] [7]), 
         .C(\register_addr[0] ), .Z(n4894[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_7_i1_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_324_4_lut (.A(n32448), .B(n32460), .C(n32511), .D(rw), 
         .Z(n32418)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_3_lut_rep_324_4_lut.init = 16'h0010;
    LUT4 i2_3_lut_3_lut_4_lut (.A(n32448), .B(n32460), .C(n32511), .D(n34320), 
         .Z(n8052)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i2_3_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i24707_2_lut_rep_298_4_lut (.A(rw), .B(n32511), .C(n32440), .D(\register_addr[0] ), 
         .Z(n32392)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i24707_2_lut_rep_298_4_lut.init = 16'h0004;
    LUT4 mux_1586_Mux_0_i1_3_lut (.A(\register[0] [0]), .B(\register[1] [0]), 
         .C(\register_addr[0] ), .Z(n4894[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(84[7] 100[14])
    defparam mux_1586_Mux_0_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_417 (.A(\select[2] ), .B(prev_select), .Z(n32511)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(82[8:29])
    defparam i1_2_lut_rep_417.init = 16'h2222;
    LUT4 i1_2_lut_2_lut_3_lut (.A(\select[2] ), .B(prev_select), .C(n34320), 
         .Z(n12099)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(82[8:29])
    defparam i1_2_lut_2_lut_3_lut.init = 16'h0202;
    FD1P3IX read_value__i0 (.D(n4894[0]), .SP(n12099), .CD(n8052), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=16, LSE_RCOL=40, LSE_LLINE=512, LSE_RLINE=522 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(73[9] 111[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i24700_2_lut_3_lut (.A(\register_addr[0] ), .B(n32418), .C(n34320), 
         .Z(n20489)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(103[9] 108[16])
    defparam i24700_2_lut_3_lut.init = 16'hf4f4;
    LUT4 i1_2_lut_3_lut (.A(\register_addr[0] ), .B(n32418), .C(n34320), 
         .Z(n12566)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(103[9] 108[16])
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i16_2_lut (.A(\select[2] ), .B(n34317), .Z(n64)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(68[19:32])
    defparam i16_2_lut.init = 16'h8888;
    PWMGenerator right (.count({Open_32, Open_33, Open_34, Open_35, 
            \count[8] , \count[7] , \count[6] , \count[5] , \count[4] , 
            \count[3] , \count[2] , \count[1] , \count[0] }), .debug_c_c(debug_c_c), 
            .n32341(n32341), .motor_pwm_r_c(motor_pwm_r_c), .GND_net(GND_net), 
            .n9633(n9633), .n14322(n14322), .\register[1] ({\register[1] }), 
            .n34320(n34320), .n3589(n3589), .n7893({n7893}), .n7902(n7902)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(118[15] 121[34])
    PWMGenerator_U6 left (.debug_c_c(debug_c_c), .n10513(n10513), .n14473(n14473), 
            .\register[0] ({\register[0] }), .count({\count[12] , \count[11] , 
            Open_36, Open_37, Open_38, Open_39, Open_40, Open_41, 
            Open_42, Open_43, Open_44, Open_45, \count[0]_adj_195 }), 
            .n32341(n32341), .\count[9] (\count[9] ), .\count[8] (\count[8]_adj_196 ), 
            .\count[6] (\count[6]_adj_197 ), .\count[5] (\count[5]_adj_198 ), 
            .\count[3] (\count[3]_adj_199 ), .\count[2] (\count[2]_adj_200 ), 
            .\count[1] (\count[1]_adj_201 ), .n34320(n34320), .motor_pwm_l_c(motor_pwm_l_c), 
            .GND_net(GND_net), .n28459(n28459), .n32356(n32356), .n10(n10), 
            .n12(n12), .\reset_count[6] (\reset_count[6] ), .n30456(n30456), 
            .\reset_count[4] (\reset_count[4] ), .\reset_count[5] (\reset_count[5] ), 
            .n30458(n30458), .\reset_count[12] (\reset_count[12] ), .\reset_count[11] (\reset_count[11] ), 
            .\reset_count[13] (\reset_count[13] ), .n29618(n29618), .n3586(n3586), 
            .n6(n6), .n32411(n32411), .n6_adj_194(n6_adj_202), .n8(n8), 
            .n7912(n7912), .n7906(n7906), .n7905(n7905), .n7908(n7908), 
            .n7910(n7910), .n7909(n7909), .n7911(n7911)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(114[15] 117[34])
    
endmodule
//
// Verilog Description of module PWMGenerator
//

module PWMGenerator (count, debug_c_c, n32341, motor_pwm_r_c, GND_net, 
            n9633, n14322, \register[1] , n34320, n3589, n7893, 
            n7902) /* synthesis syn_module_defined=1 */ ;
    output [12:0]count;
    input debug_c_c;
    input n32341;
    output motor_pwm_r_c;
    input GND_net;
    output n9633;
    input n14322;
    input [7:0]\register[1] ;
    input n34320;
    input n3589;
    output [7:0]n7893;
    output n7902;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n8031;
    wire [12:0]n43;
    
    wire n28511;
    wire [7:0]latched_width;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(15[12:25])
    wire [12:0]n28;
    wire [12:0]count_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    
    wire n30378, n19872, n17, n16, n32514, n30740, n30742, n30760, 
        n8, n27589, n27588, n27587, n27586, n27910, n27909, n27908, 
        n27907, n27906, n27905;
    
    FD1P3IX count__i0 (.D(n43[0]), .SP(n32341), .CD(n8031), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i0.GSR = "ENABLED";
    OFS1P3DX pwm_19 (.D(n28511), .SP(n32341), .SCLK(debug_c_c), .CD(GND_net), 
            .Q(motor_pwm_r_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam pwm_19.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i0 (.D(\register[1] [0]), .SP(n9633), .PD(n14322), 
            .CK(debug_c_c), .Q(latched_width[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i0.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i1 (.D(\register[1] [1]), .SP(n9633), .PD(n14322), 
            .CK(debug_c_c), .Q(latched_width[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i1.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n28[1]), .SP(n32341), .CD(n8031), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i1.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n28[2]), .SP(n32341), .CD(n8031), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n28[3]), .SP(n32341), .CD(n8031), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n28[4]), .SP(n32341), .CD(n8031), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n28[5]), .SP(n32341), .CD(n8031), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n28[6]), .SP(n32341), .CD(n8031), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n28[7]), .SP(n32341), .CD(n8031), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n28[8]), .SP(n32341), .CD(n8031), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n28[9]), .SP(n32341), .CD(n8031), .CK(debug_c_c), 
            .Q(count_c[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n28[10]), .SP(n32341), .CD(n8031), .CK(debug_c_c), 
            .Q(count_c[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i2 (.D(\register[1] [2]), .SP(n9633), .PD(n14322), 
            .CK(debug_c_c), .Q(latched_width[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i2.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i3 (.D(\register[1] [3]), .SP(n9633), .PD(n14322), 
            .CK(debug_c_c), .Q(latched_width[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i3.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i4 (.D(\register[1] [4]), .SP(n9633), .PD(n14322), 
            .CK(debug_c_c), .Q(latched_width[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i4.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i5 (.D(\register[1] [5]), .SP(n9633), .PD(n14322), 
            .CK(debug_c_c), .Q(latched_width[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i5.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i6 (.D(\register[1] [6]), .SP(n9633), .PD(n14322), 
            .CK(debug_c_c), .Q(latched_width[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i6.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n28[11]), .SP(n32341), .CD(n8031), .CK(debug_c_c), 
            .Q(count_c[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i11.GSR = "ENABLED";
    LUT4 i2274_4_lut (.A(n32341), .B(n30378), .C(n34320), .D(n19872), 
         .Z(n8031)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam i2274_4_lut.init = 16'ha0a8;
    LUT4 i9_4_lut (.A(n17), .B(count[5]), .C(n16), .D(n32514), .Z(n30378)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i9_4_lut.init = 16'h0080;
    FD1P3IX count__i12 (.D(n28[12]), .SP(n32341), .CD(n8031), .CK(debug_c_c), 
            .Q(count_c[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i12.GSR = "ENABLED";
    LUT4 i7_4_lut (.A(count[0]), .B(count_c[9]), .C(count_c[12]), .D(count[6]), 
         .Z(n17)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(count[7]), .B(count[8]), .C(count[3]), .D(count[1]), 
         .Z(n16)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i14140_2_lut (.A(count[4]), .B(count[2]), .Z(n19872)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14140_2_lut.init = 16'heeee;
    LUT4 i24254_2_lut_rep_420 (.A(count_c[10]), .B(count_c[11]), .Z(n32514)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24254_2_lut_rep_420.init = 16'heeee;
    LUT4 i24401_3_lut_4_lut (.A(count_c[10]), .B(count_c[11]), .C(n30740), 
         .D(n30742), .Z(n30760)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24401_3_lut_4_lut.init = 16'hfffe;
    FD1P3IX latched_width_i0_i7 (.D(\register[1] [7]), .SP(n9633), .CD(n14322), 
            .CK(debug_c_c), .Q(latched_width[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i7.GSR = "ENABLED";
    LUT4 i24736_4_lut (.A(count_c[11]), .B(n3589), .C(count_c[12]), .D(n8), 
         .Z(n28511)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i24736_4_lut.init = 16'h0001;
    LUT4 i2_2_lut (.A(count_c[9]), .B(count_c[10]), .Z(n8)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(26[9:19])
    defparam i2_2_lut.init = 16'heeee;
    CCU2D add_2161_9 (.A0(latched_width[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27589), .S0(n7893[7]), .S1(n7902));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2161_9.INIT0 = 16'h5555;
    defparam add_2161_9.INIT1 = 16'h0000;
    defparam add_2161_9.INJECT1_0 = "NO";
    defparam add_2161_9.INJECT1_1 = "NO";
    CCU2D add_2161_7 (.A0(latched_width[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27588), .COUT(n27589), .S0(n7893[5]), 
          .S1(n7893[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2161_7.INIT0 = 16'h5555;
    defparam add_2161_7.INIT1 = 16'h5555;
    defparam add_2161_7.INJECT1_0 = "NO";
    defparam add_2161_7.INJECT1_1 = "NO";
    CCU2D add_2161_5 (.A0(latched_width[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27587), .COUT(n27588), .S0(n7893[3]), 
          .S1(n7893[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2161_5.INIT0 = 16'h5555;
    defparam add_2161_5.INIT1 = 16'h5555;
    defparam add_2161_5.INJECT1_0 = "NO";
    defparam add_2161_5.INJECT1_1 = "NO";
    CCU2D add_2161_3 (.A0(latched_width[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27586), .COUT(n27587), .S0(n7893[1]), 
          .S1(n7893[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2161_3.INIT0 = 16'h5555;
    defparam add_2161_3.INIT1 = 16'h5555;
    defparam add_2161_3.INJECT1_0 = "NO";
    defparam add_2161_3.INJECT1_1 = "NO";
    CCU2D add_2161_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(latched_width[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27586), .S1(n7893[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2161_1.INIT0 = 16'hF000;
    defparam add_2161_1.INIT1 = 16'h5555;
    defparam add_2161_1.INJECT1_0 = "NO";
    defparam add_2161_1.INJECT1_1 = "NO";
    LUT4 i4_4_lut (.A(n30760), .B(n32341), .C(n19872), .D(count[0]), 
         .Z(n9633)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i4_4_lut.init = 16'h0004;
    LUT4 i24383_4_lut (.A(count_c[9]), .B(count[6]), .C(count[3]), .D(count[8]), 
         .Z(n30742)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24383_4_lut.init = 16'hfffe;
    LUT4 i24381_4_lut (.A(count[7]), .B(count[5]), .C(count[1]), .D(count_c[12]), 
         .Z(n30740)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24381_4_lut.init = 16'hfffe;
    CCU2D add_9_13 (.A0(count_c[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27910), .S0(n28[11]), .S1(n28[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_13.INIT0 = 16'h5aaa;
    defparam add_9_13.INIT1 = 16'h5aaa;
    defparam add_9_13.INJECT1_0 = "NO";
    defparam add_9_13.INJECT1_1 = "NO";
    CCU2D add_9_11 (.A0(count_c[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27909), .COUT(n27910), .S0(n28[9]), .S1(n28[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_11.INIT0 = 16'h5aaa;
    defparam add_9_11.INIT1 = 16'h5aaa;
    defparam add_9_11.INJECT1_0 = "NO";
    defparam add_9_11.INJECT1_1 = "NO";
    CCU2D add_9_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27908), 
          .COUT(n27909), .S0(n28[7]), .S1(n28[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_9.INIT0 = 16'h5aaa;
    defparam add_9_9.INIT1 = 16'h5aaa;
    defparam add_9_9.INJECT1_0 = "NO";
    defparam add_9_9.INJECT1_1 = "NO";
    CCU2D add_9_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27907), 
          .COUT(n27908), .S0(n28[5]), .S1(n28[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_7.INIT0 = 16'h5aaa;
    defparam add_9_7.INIT1 = 16'h5aaa;
    defparam add_9_7.INJECT1_0 = "NO";
    defparam add_9_7.INJECT1_1 = "NO";
    CCU2D add_9_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27906), 
          .COUT(n27907), .S0(n28[3]), .S1(n28[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_5.INIT0 = 16'h5aaa;
    defparam add_9_5.INIT1 = 16'h5aaa;
    defparam add_9_5.INJECT1_0 = "NO";
    defparam add_9_5.INJECT1_1 = "NO";
    CCU2D add_9_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27905), 
          .COUT(n27906), .S0(n28[1]), .S1(n28[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_3.INIT0 = 16'h5aaa;
    defparam add_9_3.INIT1 = 16'h5aaa;
    defparam add_9_3.INJECT1_0 = "NO";
    defparam add_9_3.INJECT1_1 = "NO";
    CCU2D add_9_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27905), 
          .S1(n43[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_1.INIT0 = 16'hF000;
    defparam add_9_1.INIT1 = 16'h5555;
    defparam add_9_1.INJECT1_0 = "NO";
    defparam add_9_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMGenerator_U6
//

module PWMGenerator_U6 (debug_c_c, n10513, n14473, \register[0] , count, 
            n32341, \count[9] , \count[8] , \count[6] , \count[5] , 
            \count[3] , \count[2] , \count[1] , n34320, motor_pwm_l_c, 
            GND_net, n28459, n32356, n10, n12, \reset_count[6] , 
            n30456, \reset_count[4] , \reset_count[5] , n30458, \reset_count[12] , 
            \reset_count[11] , \reset_count[13] , n29618, n3586, n6, 
            n32411, n6_adj_194, n8, n7912, n7906, n7905, n7908, 
            n7910, n7909, n7911) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    output n10513;
    input n14473;
    input [7:0]\register[0] ;
    output [12:0]count;
    input n32341;
    output \count[9] ;
    output \count[8] ;
    output \count[6] ;
    output \count[5] ;
    output \count[3] ;
    output \count[2] ;
    output \count[1] ;
    input n34320;
    output motor_pwm_l_c;
    input GND_net;
    input n28459;
    output n32356;
    input n10;
    output n12;
    input \reset_count[6] ;
    input n30456;
    input \reset_count[4] ;
    input \reset_count[5] ;
    output n30458;
    input \reset_count[12] ;
    input \reset_count[11] ;
    input \reset_count[13] ;
    output n29618;
    input n3586;
    output n6;
    output n32411;
    input n6_adj_194;
    output n8;
    output n7912;
    output n7906;
    output n7905;
    output n7908;
    output n7910;
    output n7909;
    output n7911;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [7:0]latched_width;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(15[12:25])
    wire [12:0]n42;
    
    wire n8027;
    wire [12:0]n43;
    wire [12:0]count_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    wire [12:0]n28;
    
    wire n28537, n30611, n15_adj_384, n14, n32492, n30724, n30752;
    wire [7:0]n7903;
    
    wire n30728, n27903, n27902, n27901, n27900, n27899, n27898, 
        n27897, n27896, n27895, n27894;
    
    FD1P3JX latched_width_i0_i2 (.D(\register[0] [2]), .SP(n10513), .PD(n14473), 
            .CK(debug_c_c), .Q(latched_width[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i2.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i1 (.D(\register[0] [1]), .SP(n10513), .PD(n14473), 
            .CK(debug_c_c), .Q(latched_width[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i1.GSR = "ENABLED";
    FD1P3AX count__i0 (.D(n42[0]), .SP(n32341), .CK(debug_c_c), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i0.GSR = "ENABLED";
    FD1P3IX count__i12 (.D(n43[12]), .SP(n32341), .CD(n8027), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i12.GSR = "ENABLED";
    FD1P3IX count__i11 (.D(n43[11]), .SP(n32341), .CD(n8027), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i11.GSR = "ENABLED";
    FD1P3IX count__i10 (.D(n43[10]), .SP(n32341), .CD(n8027), .CK(debug_c_c), 
            .Q(count_c[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i10.GSR = "ENABLED";
    FD1P3IX count__i9 (.D(n43[9]), .SP(n32341), .CD(n8027), .CK(debug_c_c), 
            .Q(\count[9] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i9.GSR = "ENABLED";
    FD1P3IX count__i8 (.D(n43[8]), .SP(n32341), .CD(n8027), .CK(debug_c_c), 
            .Q(\count[8] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i8.GSR = "ENABLED";
    FD1P3IX count__i7 (.D(n43[7]), .SP(n32341), .CD(n8027), .CK(debug_c_c), 
            .Q(count_c[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i7.GSR = "ENABLED";
    FD1P3IX count__i6 (.D(n43[6]), .SP(n32341), .CD(n8027), .CK(debug_c_c), 
            .Q(\count[6] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i6.GSR = "ENABLED";
    FD1P3IX count__i5 (.D(n43[5]), .SP(n32341), .CD(n8027), .CK(debug_c_c), 
            .Q(\count[5] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i5.GSR = "ENABLED";
    FD1P3IX count__i4 (.D(n43[4]), .SP(n32341), .CD(n8027), .CK(debug_c_c), 
            .Q(count_c[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i4.GSR = "ENABLED";
    FD1P3IX count__i3 (.D(n43[3]), .SP(n32341), .CD(n8027), .CK(debug_c_c), 
            .Q(\count[3] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i3.GSR = "ENABLED";
    FD1P3IX count__i2 (.D(n43[2]), .SP(n32341), .CD(n8027), .CK(debug_c_c), 
            .Q(\count[2] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i2.GSR = "ENABLED";
    FD1P3IX count__i1 (.D(n43[1]), .SP(n32341), .CD(n8027), .CK(debug_c_c), 
            .Q(\count[1] ));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam count__i1.GSR = "ENABLED";
    LUT4 i14007_2_lut (.A(n28[0]), .B(n8027), .Z(n42[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam i14007_2_lut.init = 16'h2222;
    LUT4 i2270_4_lut (.A(n32341), .B(n28537), .C(n34320), .D(n30611), 
         .Z(n8027)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam i2270_4_lut.init = 16'ha0a8;
    LUT4 i8_4_lut (.A(n15_adj_384), .B(\count[8] ), .C(n14), .D(\count[9] ), 
         .Z(n28537)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(\count[5] ), .B(\count[6] ), .C(count[0]), .D(\count[1] ), 
         .Z(n15_adj_384)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_3_lut (.A(count[12]), .B(count_c[7]), .C(\count[3] ), .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5_3_lut.init = 16'h8080;
    LUT4 i2_4_lut (.A(n32341), .B(n32492), .C(n30724), .D(n30752), .Z(n10513)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i2_4_lut.init = 16'h0002;
    FD1P3JX latched_width_i0_i0 (.D(\register[0] [0]), .SP(n10513), .PD(n14473), 
            .CK(debug_c_c), .Q(latched_width[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i0.GSR = "ENABLED";
    FD1P3IX pwm_19 (.D(n28459), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(motor_pwm_l_c));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam pwm_19.GSR = "ENABLED";
    LUT4 i10_2_lut_rep_262 (.A(n7903[7]), .B(count_c[7]), .Z(n32356)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    defparam i10_2_lut_rep_262.init = 16'h6666;
    LUT4 LessThan_1434_i12_3_lut_3_lut (.A(n7903[7]), .B(count_c[7]), .C(n10), 
         .Z(n12)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    defparam LessThan_1434_i12_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i45_2_lut_rep_398 (.A(\count[2] ), .B(count_c[4]), .Z(n32492)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i45_2_lut_rep_398.init = 16'heeee;
    LUT4 i24256_3_lut_4_lut (.A(\count[2] ), .B(count_c[4]), .C(count[11]), 
         .D(count_c[10]), .Z(n30611)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24256_3_lut_4_lut.init = 16'hfffe;
    LUT4 i24365_4_lut (.A(count[11]), .B(count_c[7]), .C(\count[5] ), 
         .D(\count[9] ), .Z(n30724)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24365_4_lut.init = 16'hfffe;
    LUT4 i24393_4_lut (.A(count[12]), .B(n30728), .C(\count[8] ), .D(count[0]), 
         .Z(n30752)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24393_4_lut.init = 16'hfffe;
    LUT4 i24369_4_lut (.A(\count[3] ), .B(count_c[10]), .C(\count[1] ), 
         .D(\count[6] ), .Z(n30728)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24369_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut (.A(\reset_count[6] ), .B(n30456), .C(\reset_count[4] ), 
         .D(\reset_count[5] ), .Z(n30458)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'heeec;
    LUT4 i2_3_lut (.A(\reset_count[12] ), .B(\reset_count[11] ), .C(\reset_count[13] ), 
         .Z(n29618)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut (.A(count_c[10]), .B(n3586), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(26[9:19])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i9_2_lut_rep_317 (.A(n7903[4]), .B(count_c[4]), .Z(n32411)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    defparam i9_2_lut_rep_317.init = 16'h6666;
    LUT4 LessThan_1434_i8_3_lut_3_lut (.A(n7903[4]), .B(count_c[4]), .C(n6_adj_194), 
         .Z(n8)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(14[13:18])
    defparam LessThan_1434_i8_3_lut_3_lut.init = 16'hd4d4;
    FD1P3IX latched_width_i0_i7 (.D(\register[0] [7]), .SP(n10513), .CD(n14473), 
            .CK(debug_c_c), .Q(latched_width[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i7.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i6 (.D(\register[0] [6]), .SP(n10513), .PD(n14473), 
            .CK(debug_c_c), .Q(latched_width[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i6.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i5 (.D(\register[0] [5]), .SP(n10513), .PD(n14473), 
            .CK(debug_c_c), .Q(latched_width[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i5.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i4 (.D(\register[0] [4]), .SP(n10513), .PD(n14473), 
            .CK(debug_c_c), .Q(latched_width[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i4.GSR = "ENABLED";
    FD1P3JX latched_width_i0_i3 (.D(\register[0] [3]), .SP(n10513), .PD(n14473), 
            .CK(debug_c_c), .Q(latched_width[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(17[9] 38[6])
    defparam latched_width_i0_i3.GSR = "ENABLED";
    CCU2D add_9_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27903), .S0(n43[11]), .S1(n43[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_13.INIT0 = 16'h5aaa;
    defparam add_9_13.INIT1 = 16'h5aaa;
    defparam add_9_13.INJECT1_0 = "NO";
    defparam add_9_13.INJECT1_1 = "NO";
    CCU2D add_9_11 (.A0(\count[9] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27902), .COUT(n27903), .S0(n43[9]), .S1(n43[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_11.INIT0 = 16'h5aaa;
    defparam add_9_11.INIT1 = 16'h5aaa;
    defparam add_9_11.INJECT1_0 = "NO";
    defparam add_9_11.INJECT1_1 = "NO";
    CCU2D add_9_9 (.A0(count_c[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count[8] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27901), .COUT(n27902), .S0(n43[7]), .S1(n43[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_9.INIT0 = 16'h5aaa;
    defparam add_9_9.INIT1 = 16'h5aaa;
    defparam add_9_9.INJECT1_0 = "NO";
    defparam add_9_9.INJECT1_1 = "NO";
    CCU2D add_9_7 (.A0(\count[5] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count[6] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27900), .COUT(n27901), .S0(n43[5]), .S1(n43[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_7.INIT0 = 16'h5aaa;
    defparam add_9_7.INIT1 = 16'h5aaa;
    defparam add_9_7.INJECT1_0 = "NO";
    defparam add_9_7.INJECT1_1 = "NO";
    CCU2D add_9_5 (.A0(\count[3] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_c[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27899), .COUT(n27900), .S0(n43[3]), .S1(n43[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_5.INIT0 = 16'h5aaa;
    defparam add_9_5.INIT1 = 16'h5aaa;
    defparam add_9_5.INJECT1_0 = "NO";
    defparam add_9_5.INJECT1_1 = "NO";
    CCU2D add_9_3 (.A0(\count[1] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count[2] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27898), .COUT(n27899), .S0(n43[1]), .S1(n43[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_3.INIT0 = 16'h5aaa;
    defparam add_9_3.INIT1 = 16'h5aaa;
    defparam add_9_3.INJECT1_0 = "NO";
    defparam add_9_3.INJECT1_1 = "NO";
    CCU2D add_9_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27898), 
          .S1(n28[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(36[16:25])
    defparam add_9_1.INIT0 = 16'hF000;
    defparam add_9_1.INIT1 = 16'h5555;
    defparam add_9_1.INJECT1_0 = "NO";
    defparam add_9_1.INJECT1_1 = "NO";
    CCU2D add_2162_9 (.A0(latched_width[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27897), .S0(n7903[7]), .S1(n7912));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2162_9.INIT0 = 16'h5555;
    defparam add_2162_9.INIT1 = 16'h0000;
    defparam add_2162_9.INJECT1_0 = "NO";
    defparam add_2162_9.INJECT1_1 = "NO";
    CCU2D add_2162_7 (.A0(latched_width[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27896), .COUT(n27897), .S0(n7906), .S1(n7905));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2162_7.INIT0 = 16'h5555;
    defparam add_2162_7.INIT1 = 16'h5555;
    defparam add_2162_7.INJECT1_0 = "NO";
    defparam add_2162_7.INJECT1_1 = "NO";
    CCU2D add_2162_5 (.A0(latched_width[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27895), .COUT(n27896), .S0(n7908), .S1(n7903[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2162_5.INIT0 = 16'h5555;
    defparam add_2162_5.INIT1 = 16'h5555;
    defparam add_2162_5.INJECT1_0 = "NO";
    defparam add_2162_5.INJECT1_1 = "NO";
    CCU2D add_2162_3 (.A0(latched_width[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(latched_width[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27894), .COUT(n27895), .S0(n7910), .S1(n7909));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2162_3.INIT0 = 16'h5555;
    defparam add_2162_3.INIT1 = 16'h5555;
    defparam add_2162_3.INJECT1_0 = "NO";
    defparam add_2162_3.INJECT1_1 = "NO";
    CCU2D add_2162_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(latched_width[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27894), .S1(n7911));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(28[18:43])
    defparam add_2162_1.INIT0 = 16'hF000;
    defparam add_2162_1.INIT1 = 16'h5555;
    defparam add_2162_1.INJECT1_0 = "NO";
    defparam add_2162_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module GlobalControlPeripheral
//

module GlobalControlPeripheral (n32448, n32504, n11645, register_addr, 
            read_value, debug_c_c, n32379, n11753, n30258, n8048, 
            n21, n15, read_size, n302, \register[2][0] , n34321, 
            \register[0][2] , \select[1] , n34323, n34322, \register[2][3] , 
            n28356, n32422, n32433, n32429, n4, n34317, n32472, 
            rw, n6, force_pause, \databus[1] , n34320, n20268, xbee_pause_c, 
            n10513, n14473, signal_light_c, \control_reg[7] , n28309, 
            stepping, n9633, n14322, \control_reg[7]_adj_188 , n28270, 
            stepping_adj_189, \control_reg[7]_adj_190 , n28332, n21_adj_191, 
            \control_reg[7]_adj_192 , n28296, stepping_adj_193, n32503, 
            n32455, \select[4] , n32439, n32443, GND_net) /* synthesis syn_module_defined=1 */ ;
    input n32448;
    input n32504;
    input n11645;
    input [7:0]register_addr;
    output [31:0]read_value;
    input debug_c_c;
    output n32379;
    input n11753;
    output n30258;
    input n8048;
    input n21;
    input n15;
    output [2:0]read_size;
    input n302;
    output \register[2][0] ;
    input n34321;
    output \register[0][2] ;
    input \select[1] ;
    input n34323;
    input n34322;
    output \register[2][3] ;
    input n28356;
    input n32422;
    input n32433;
    input n32429;
    input n4;
    input n34317;
    output n32472;
    input rw;
    output n6;
    output force_pause;
    input \databus[1] ;
    input n34320;
    output n20268;
    input xbee_pause_c;
    input n10513;
    output n14473;
    output signal_light_c;
    input \control_reg[7] ;
    input n28309;
    output stepping;
    input n9633;
    output n14322;
    input \control_reg[7]_adj_188 ;
    input n28270;
    output stepping_adj_189;
    input \control_reg[7]_adj_190 ;
    input n28332;
    output n21_adj_191;
    input \control_reg[7]_adj_192 ;
    input n28296;
    output stepping_adj_193;
    output n32503;
    output n32455;
    input \select[4] ;
    output n32439;
    input n32443;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(23[14:22])
    
    wire n29649, n29638, n29637, n29635, n29650, n29628, n29631, 
        n29654, n29629, n30168, n29647, n29646, n29644, n29639, 
        n29651, n29632, n29634, n30418, n29630, n29642, n29645, 
        n29641, n29633, n29655, n29640, n29652, n29636, n29653, 
        n29648, n29643, n30417, n32334;
    wire [31:0]read_value_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(30[13:23])
    
    wire n32335, n24, n7999;
    wire [31:0]n100;
    
    wire prev_clk_1Hz, clk_1Hz, n178, prev_select, n32512, n14414, 
        n14413, n32485, n27997, n32479, n27, n27_adj_376, n16, 
        n16_adj_383, n27569, n27568, n27567, n27566, n27565, n27564, 
        n27563, n27562, n27561, n27560, n27559, n27558, n27557, 
        n27556, n27555, n27554;
    
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32448), .B(n32504), .C(\register[2] [19]), 
         .D(n11645), .Z(n29649)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_436 (.A(n32448), .B(n32504), .C(\register[2] [20]), 
         .D(n11645), .Z(n29638)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_436.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_437 (.A(n32448), .B(n32504), .C(\register[2] [29]), 
         .D(n11645), .Z(n29637)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_437.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_438 (.A(n32448), .B(n32504), .C(\register[2] [21]), 
         .D(n11645), .Z(n29635)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_438.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_439 (.A(n32448), .B(n32504), .C(\register[2] [22]), 
         .D(n11645), .Z(n29650)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_439.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_440 (.A(n32448), .B(n32504), .C(\register[2] [23]), 
         .D(n11645), .Z(n29628)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_440.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_441 (.A(n32448), .B(n32504), .C(\register[2] [24]), 
         .D(n11645), .Z(n29631)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_441.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_442 (.A(n32448), .B(n32504), .C(\register[2] [25]), 
         .D(n11645), .Z(n29654)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_442.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_443 (.A(n32448), .B(n32504), .C(\register[2] [26]), 
         .D(n11645), .Z(n29629)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_443.init = 16'h1000;
    LUT4 i1_3_lut_4_lut (.A(n32448), .B(n32504), .C(register_addr[0]), 
         .D(register_addr[1]), .Z(n30168)) /* synthesis lut_function=(!(A+(B+!((D)+!C)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h1101;
    LUT4 i1_2_lut_3_lut_4_lut_adj_444 (.A(n32448), .B(n32504), .C(\register[2] [30]), 
         .D(n11645), .Z(n29647)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_444.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_445 (.A(n32448), .B(n32504), .C(\register[2] [31]), 
         .D(n11645), .Z(n29646)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_445.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_446 (.A(n32448), .B(n32504), .C(\register[2] [28]), 
         .D(n11645), .Z(n29644)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_446.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_447 (.A(n32448), .B(n32504), .C(\register[2] [5]), 
         .D(n11645), .Z(n29639)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_447.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_448 (.A(n32448), .B(n32504), .C(\register[2] [7]), 
         .D(n11645), .Z(n29651)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_448.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_449 (.A(n32448), .B(n32504), .C(\register[2] [16]), 
         .D(n11645), .Z(n29632)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_449.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_450 (.A(n32448), .B(n32504), .C(\register[2] [27]), 
         .D(n11645), .Z(n29634)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_450.init = 16'h1000;
    FD1P3AX read_value__i0 (.D(n30418), .SP(n32379), .CK(debug_c_c), .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(n11753), .B(register_addr[3]), .Z(n30258)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam i1_2_lut.init = 16'h2222;
    FD1P3IX read_value__i31 (.D(n29646), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX read_value__i30 (.D(n29647), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3IX read_value__i29 (.D(n29637), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3IX read_value__i28 (.D(n29644), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3IX read_value__i27 (.D(n29634), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3IX read_value__i26 (.D(n29629), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3IX read_value__i25 (.D(n29654), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3IX read_value__i24 (.D(n29631), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3IX read_value__i23 (.D(n29628), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3IX read_value__i22 (.D(n29650), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3IX read_value__i21 (.D(n29635), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3IX read_value__i20 (.D(n29638), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3IX read_value__i19 (.D(n29649), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3IX read_value__i18 (.D(n29630), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n29642), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n29632), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n29645), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3IX read_value__i14 (.D(n29641), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3IX read_value__i13 (.D(n29633), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3IX read_value__i12 (.D(n29655), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3IX read_value__i11 (.D(n29640), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3IX read_value__i10 (.D(n29652), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3IX read_value__i9 (.D(n29636), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3IX read_value__i8 (.D(n29653), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n29651), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n29648), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n29639), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n29643), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n30417), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n32334), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n32335), .SP(n32379), .CD(n8048), .CK(debug_c_c), 
            .Q(read_value_c[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_value__i1.GSR = "ENABLED";
    PFUMX i33 (.BLUT(n21), .ALUT(n15), .C0(register_addr[1]), .Z(n24));
    FD1P3AX read_size_i0_i0 (.D(n302), .SP(n32379), .CK(debug_c_c), .Q(read_size[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i0.GSR = "ENABLED";
    FD1P3IX uptime_count__i0 (.D(n100[0]), .SP(n7999), .CD(n34321), .CK(debug_c_c), 
            .Q(\register[2][0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i0.GSR = "ENABLED";
    FD1S3AX prev_clk_1Hz_149 (.D(clk_1Hz), .CK(debug_c_c), .Q(prev_clk_1Hz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam prev_clk_1Hz_149.GSR = "ENABLED";
    FD1S3AX xbee_pause_latched_150 (.D(n178), .CK(debug_c_c), .Q(\register[0][2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam xbee_pause_latched_150.GSR = "ENABLED";
    FD1S3AX prev_select_148 (.D(\select[1] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam prev_select_148.GSR = "ENABLED";
    FD1P3IX uptime_count__i31 (.D(n100[31]), .SP(n7999), .CD(n34323), 
            .CK(debug_c_c), .Q(\register[2] [31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i31.GSR = "ENABLED";
    FD1P3IX uptime_count__i30 (.D(n100[30]), .SP(n7999), .CD(n34321), 
            .CK(debug_c_c), .Q(\register[2] [30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i30.GSR = "ENABLED";
    FD1P3IX uptime_count__i29 (.D(n100[29]), .SP(n7999), .CD(n34321), 
            .CK(debug_c_c), .Q(\register[2] [29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i29.GSR = "ENABLED";
    FD1P3IX uptime_count__i28 (.D(n100[28]), .SP(n7999), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i28.GSR = "ENABLED";
    FD1P3IX uptime_count__i27 (.D(n100[27]), .SP(n7999), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i27.GSR = "ENABLED";
    FD1P3IX uptime_count__i26 (.D(n100[26]), .SP(n7999), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i26.GSR = "ENABLED";
    FD1P3IX uptime_count__i25 (.D(n100[25]), .SP(n7999), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i25.GSR = "ENABLED";
    FD1P3IX uptime_count__i24 (.D(n100[24]), .SP(n7999), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i24.GSR = "ENABLED";
    FD1P3IX uptime_count__i23 (.D(n100[23]), .SP(n7999), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i23.GSR = "ENABLED";
    FD1P3IX uptime_count__i22 (.D(n100[22]), .SP(n7999), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i22.GSR = "ENABLED";
    FD1P3IX uptime_count__i21 (.D(n100[21]), .SP(n7999), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i21.GSR = "ENABLED";
    FD1P3IX uptime_count__i20 (.D(n100[20]), .SP(n7999), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i20.GSR = "ENABLED";
    FD1P3IX uptime_count__i19 (.D(n100[19]), .SP(n7999), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i19.GSR = "ENABLED";
    FD1P3IX uptime_count__i18 (.D(n100[18]), .SP(n7999), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i18.GSR = "ENABLED";
    FD1P3IX uptime_count__i17 (.D(n100[17]), .SP(n7999), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i17.GSR = "ENABLED";
    FD1P3IX uptime_count__i16 (.D(n100[16]), .SP(n7999), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i16.GSR = "ENABLED";
    FD1P3IX uptime_count__i15 (.D(n100[15]), .SP(n7999), .CD(n34321), 
            .CK(debug_c_c), .Q(\register[2] [15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i15.GSR = "ENABLED";
    FD1P3IX uptime_count__i14 (.D(n100[14]), .SP(n7999), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i14.GSR = "ENABLED";
    FD1P3IX uptime_count__i13 (.D(n100[13]), .SP(n7999), .CD(n34321), 
            .CK(debug_c_c), .Q(\register[2] [13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i13.GSR = "ENABLED";
    FD1P3IX uptime_count__i12 (.D(n100[12]), .SP(n32512), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i12.GSR = "ENABLED";
    FD1P3IX uptime_count__i11 (.D(n100[11]), .SP(n7999), .CD(n34322), 
            .CK(debug_c_c), .Q(\register[2] [11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i11.GSR = "ENABLED";
    FD1P3IX uptime_count__i10 (.D(n100[10]), .SP(n7999), .CD(n34321), 
            .CK(debug_c_c), .Q(\register[2] [10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i10.GSR = "ENABLED";
    FD1P3IX uptime_count__i9 (.D(n100[9]), .SP(n7999), .CD(n34322), .CK(debug_c_c), 
            .Q(\register[2] [9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i9.GSR = "ENABLED";
    FD1P3IX uptime_count__i8 (.D(n100[8]), .SP(n7999), .CD(n34321), .CK(debug_c_c), 
            .Q(\register[2] [8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i8.GSR = "ENABLED";
    FD1P3IX uptime_count__i7 (.D(n100[7]), .SP(n7999), .CD(n34322), .CK(debug_c_c), 
            .Q(\register[2] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i7.GSR = "ENABLED";
    FD1P3IX uptime_count__i6 (.D(n100[6]), .SP(n7999), .CD(n34322), .CK(debug_c_c), 
            .Q(\register[2] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i6.GSR = "ENABLED";
    FD1P3IX uptime_count__i5 (.D(n100[5]), .SP(n7999), .CD(n34322), .CK(debug_c_c), 
            .Q(\register[2] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i5.GSR = "ENABLED";
    FD1P3IX uptime_count__i4 (.D(n100[4]), .SP(n7999), .CD(n34322), .CK(debug_c_c), 
            .Q(\register[2] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i4.GSR = "ENABLED";
    FD1P3IX uptime_count__i3 (.D(n100[3]), .SP(n7999), .CD(n34321), .CK(debug_c_c), 
            .Q(\register[2][3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i3.GSR = "ENABLED";
    FD1P3IX read_size_i0_i1 (.D(n28356), .SP(n32379), .CD(n14414), .CK(debug_c_c), 
            .Q(read_size[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i1.GSR = "ENABLED";
    FD1P3IX read_size_i0_i2 (.D(n32422), .SP(n32379), .CD(n14413), .CK(debug_c_c), 
            .Q(read_size[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam read_size_i0_i2.GSR = "ENABLED";
    FD1P3IX uptime_count__i2 (.D(n100[2]), .SP(n7999), .CD(n32433), .CK(debug_c_c), 
            .Q(\register[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i2.GSR = "ENABLED";
    FD1P3IX uptime_count__i1 (.D(n100[1]), .SP(n7999), .CD(n32433), .CK(debug_c_c), 
            .Q(\register[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=45, LSE_RCOL=74, LSE_LLINE=495, LSE_RLINE=505 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam uptime_count__i1.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n32485), .B(n32429), .C(n4), .D(register_addr[1]), 
         .Z(n30417)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h3011;
    LUT4 i14_2_lut_rep_378 (.A(\select[1] ), .B(n34317), .Z(n32472)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(35[19:32])
    defparam i14_2_lut_rep_378.init = 16'h8888;
    LUT4 Select_3624_i6_2_lut_3_lut (.A(\select[1] ), .B(rw), .C(read_value_c[1]), 
         .Z(n6)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(35[19:32])
    defparam Select_3624_i6_2_lut_3_lut.init = 16'h8080;
    FD1P3IX force_pause_151 (.D(\databus[1] ), .SP(n27997), .CD(n32433), 
            .CK(debug_c_c), .Q(force_pause));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam force_pause_151.GSR = "ENABLED";
    LUT4 i117_2_lut_rep_385 (.A(prev_select), .B(\select[1] ), .Z(n32479)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(62[9:30])
    defparam i117_2_lut_rep_385.init = 16'h4444;
    LUT4 i8648_2_lut_3_lut_3_lut_4_lut (.A(prev_select), .B(\select[1] ), 
         .C(n30168), .D(n34320), .Z(n14414)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(62[9:30])
    defparam i8648_2_lut_3_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i8647_2_lut_3_lut_3_lut_4_lut (.A(prev_select), .B(\select[1] ), 
         .C(n30168), .D(n34320), .Z(n14413)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(62[9:30])
    defparam i8647_2_lut_3_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i889_2_lut_rep_285_2_lut_3_lut (.A(prev_select), .B(\select[1] ), 
         .C(n34320), .Z(n32379)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(62[9:30])
    defparam i889_2_lut_rep_285_2_lut_3_lut.init = 16'h0404;
    LUT4 i1_3_lut_4_lut_adj_451 (.A(register_addr[0]), .B(n32448), .C(n24), 
         .D(n8048), .Z(n30418)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_3_lut_4_lut_adj_451.init = 16'h0010;
    LUT4 i14532_3_lut (.A(register_addr[2]), .B(register_addr[1]), .C(register_addr[0]), 
         .Z(n20268)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i14532_3_lut.init = 16'ha8a8;
    LUT4 i24258_2_lut_rep_391 (.A(register_addr[3]), .B(register_addr[2]), 
         .Z(n32485)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i24258_2_lut_rep_391.init = 16'hbbbb;
    LUT4 i1_3_lut_4_lut_adj_452 (.A(register_addr[3]), .B(register_addr[2]), 
         .C(\register[0][2] ), .D(register_addr[0]), .Z(n27)) /* synthesis lut_function=(A (C+(D))+!A (B (D)+!B (C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_452.init = 16'hffb0;
    LUT4 i1_3_lut_4_lut_adj_453 (.A(register_addr[3]), .B(register_addr[2]), 
         .C(force_pause), .D(register_addr[0]), .Z(n27_adj_376)) /* synthesis lut_function=(A (C+(D))+!A (B (D)+!B (C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_453.init = 16'hffb0;
    LUT4 i114_1_lut (.A(xbee_pause_c), .Z(n178)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(54[26:39])
    defparam i114_1_lut.init = 16'h5555;
    LUT4 i8712_2_lut_3_lut (.A(\register[0][2] ), .B(force_pause), .C(n10513), 
         .Z(n14473)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i8712_2_lut_3_lut.init = 16'he0e0;
    LUT4 i13928_2_lut_3_lut (.A(\register[0][2] ), .B(force_pause), .C(clk_1Hz), 
         .Z(signal_light_c)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i13928_2_lut_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_4_lut (.A(\register[0][2] ), .B(force_pause), .C(\control_reg[7] ), 
         .D(n28309), .Z(stepping)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut.init = 16'h1000;
    LUT4 i8679_2_lut_3_lut (.A(\register[0][2] ), .B(force_pause), .C(n9633), 
         .Z(n14322)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i8679_2_lut_3_lut.init = 16'he0e0;
    LUT4 i2_3_lut_4_lut_adj_454 (.A(\register[0][2] ), .B(force_pause), 
         .C(\control_reg[7]_adj_188 ), .D(n28270), .Z(stepping_adj_189)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_454.init = 16'h1000;
    LUT4 i2_3_lut_4_lut_adj_455 (.A(\register[0][2] ), .B(force_pause), 
         .C(\control_reg[7]_adj_190 ), .D(n28332), .Z(n21_adj_191)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_455.init = 16'h1000;
    LUT4 i2_3_lut_4_lut_adj_456 (.A(\register[0][2] ), .B(force_pause), 
         .C(\control_reg[7]_adj_192 ), .D(n28296), .Z(stepping_adj_193)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(38[24:56])
    defparam i2_3_lut_4_lut_adj_456.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_457 (.A(n32448), .B(n32504), .C(\register[2] [6]), 
         .D(n11645), .Z(n29648)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_457.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_458 (.A(n32448), .B(n32504), .C(\register[2] [4]), 
         .D(n11645), .Z(n29643)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_458.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_459 (.A(n32448), .B(n32504), .C(\register[2] [8]), 
         .D(n11645), .Z(n29653)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_459.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_460 (.A(n32448), .B(n32504), .C(\register[2] [9]), 
         .D(n11645), .Z(n29636)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_460.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_461 (.A(n32448), .B(n32504), .C(\register[2] [10]), 
         .D(n11645), .Z(n29652)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_461.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_462 (.A(n32448), .B(n32504), .C(\register[2] [11]), 
         .D(n11645), .Z(n29640)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_462.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_463 (.A(n32448), .B(n32504), .C(\register[2] [12]), 
         .D(n11645), .Z(n29655)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_463.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_464 (.A(n32448), .B(n32504), .C(\register[2] [13]), 
         .D(n11645), .Z(n29633)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_464.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_465 (.A(n32448), .B(n32504), .C(\register[2] [14]), 
         .D(n11645), .Z(n29641)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_465.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_466 (.A(n32448), .B(n32504), .C(\register[2] [15]), 
         .D(n11645), .Z(n29645)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_466.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_467 (.A(n32448), .B(n32504), .C(\register[2] [17]), 
         .D(n11645), .Z(n29642)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_467.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_468 (.A(n32448), .B(n32504), .C(\register[2] [18]), 
         .D(n11645), .Z(n29630)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_468.init = 16'h1000;
    LUT4 i13813_2_lut_rep_409 (.A(register_addr[7]), .B(register_addr[6]), 
         .Z(n32503)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13813_2_lut_rep_409.init = 16'heeee;
    LUT4 i1_2_lut_rep_361_3_lut_4_lut (.A(register_addr[7]), .B(register_addr[6]), 
         .C(register_addr[5]), .D(register_addr[4]), .Z(n32455)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_361_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_345_3_lut_4_lut (.A(register_addr[7]), .B(register_addr[6]), 
         .C(\select[4] ), .D(n32504), .Z(n32439)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_345_3_lut_4_lut.init = 16'h0010;
    LUT4 i134_2_lut_rep_418 (.A(prev_clk_1Hz), .B(clk_1Hz), .Z(n32512)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(102[9:32])
    defparam i134_2_lut_rep_418.init = 16'h4444;
    LUT4 i2256_2_lut_3_lut (.A(prev_clk_1Hz), .B(clk_1Hz), .C(n34320), 
         .Z(n7999)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(102[9:32])
    defparam i2256_2_lut_3_lut.init = 16'hf4f4;
    LUT4 i2_4_lut (.A(n34320), .B(rw), .C(n32479), .D(n32422), .Z(n27997)) /* synthesis lut_function=(!(A (B+(D))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(50[9] 105[6])
    defparam i2_4_lut.init = 16'h0032;
    LUT4 n27_bdd_4_lut (.A(n27), .B(n16), .C(register_addr[1]), .D(n32443), 
         .Z(n32334)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n27_bdd_4_lut.init = 16'h00ca;
    LUT4 i1_2_lut_adj_469 (.A(\register[2] [2]), .B(register_addr[0]), .Z(n16)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_469.init = 16'h2222;
    LUT4 i1_2_lut_adj_470 (.A(\register[2] [1]), .B(register_addr[0]), .Z(n16_adj_383)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_470.init = 16'h2222;
    LUT4 n27_bdd_4_lut_adj_471 (.A(n27_adj_376), .B(n16_adj_383), .C(register_addr[1]), 
         .D(n32443), .Z(n32335)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n27_bdd_4_lut_adj_471.init = 16'h00ca;
    CCU2D add_134_33 (.A0(\register[2] [31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27569), .S0(n100[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_33.INIT0 = 16'h5aaa;
    defparam add_134_33.INIT1 = 16'h0000;
    defparam add_134_33.INJECT1_0 = "NO";
    defparam add_134_33.INJECT1_1 = "NO";
    CCU2D add_134_31 (.A0(\register[2] [29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27568), .COUT(n27569), .S0(n100[29]), 
          .S1(n100[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_31.INIT0 = 16'h5aaa;
    defparam add_134_31.INIT1 = 16'h5aaa;
    defparam add_134_31.INJECT1_0 = "NO";
    defparam add_134_31.INJECT1_1 = "NO";
    CCU2D add_134_29 (.A0(\register[2] [27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27567), .COUT(n27568), .S0(n100[27]), 
          .S1(n100[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_29.INIT0 = 16'h5aaa;
    defparam add_134_29.INIT1 = 16'h5aaa;
    defparam add_134_29.INJECT1_0 = "NO";
    defparam add_134_29.INJECT1_1 = "NO";
    CCU2D add_134_27 (.A0(\register[2] [25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27566), .COUT(n27567), .S0(n100[25]), 
          .S1(n100[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_27.INIT0 = 16'h5aaa;
    defparam add_134_27.INIT1 = 16'h5aaa;
    defparam add_134_27.INJECT1_0 = "NO";
    defparam add_134_27.INJECT1_1 = "NO";
    CCU2D add_134_25 (.A0(\register[2] [23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27565), .COUT(n27566), .S0(n100[23]), 
          .S1(n100[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_25.INIT0 = 16'h5aaa;
    defparam add_134_25.INIT1 = 16'h5aaa;
    defparam add_134_25.INJECT1_0 = "NO";
    defparam add_134_25.INJECT1_1 = "NO";
    CCU2D add_134_23 (.A0(\register[2] [21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27564), .COUT(n27565), .S0(n100[21]), 
          .S1(n100[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_23.INIT0 = 16'h5aaa;
    defparam add_134_23.INIT1 = 16'h5aaa;
    defparam add_134_23.INJECT1_0 = "NO";
    defparam add_134_23.INJECT1_1 = "NO";
    CCU2D add_134_21 (.A0(\register[2] [19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27563), .COUT(n27564), .S0(n100[19]), 
          .S1(n100[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_21.INIT0 = 16'h5aaa;
    defparam add_134_21.INIT1 = 16'h5aaa;
    defparam add_134_21.INJECT1_0 = "NO";
    defparam add_134_21.INJECT1_1 = "NO";
    CCU2D add_134_19 (.A0(\register[2] [17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27562), .COUT(n27563), .S0(n100[17]), 
          .S1(n100[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_19.INIT0 = 16'h5aaa;
    defparam add_134_19.INIT1 = 16'h5aaa;
    defparam add_134_19.INJECT1_0 = "NO";
    defparam add_134_19.INJECT1_1 = "NO";
    CCU2D add_134_17 (.A0(\register[2] [15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27561), .COUT(n27562), .S0(n100[15]), 
          .S1(n100[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_17.INIT0 = 16'h5aaa;
    defparam add_134_17.INIT1 = 16'h5aaa;
    defparam add_134_17.INJECT1_0 = "NO";
    defparam add_134_17.INJECT1_1 = "NO";
    CCU2D add_134_15 (.A0(\register[2] [13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27560), .COUT(n27561), .S0(n100[13]), 
          .S1(n100[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_15.INIT0 = 16'h5aaa;
    defparam add_134_15.INIT1 = 16'h5aaa;
    defparam add_134_15.INJECT1_0 = "NO";
    defparam add_134_15.INJECT1_1 = "NO";
    CCU2D add_134_13 (.A0(\register[2] [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27559), .COUT(n27560), .S0(n100[11]), 
          .S1(n100[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_13.INIT0 = 16'h5aaa;
    defparam add_134_13.INIT1 = 16'h5aaa;
    defparam add_134_13.INJECT1_0 = "NO";
    defparam add_134_13.INJECT1_1 = "NO";
    CCU2D add_134_11 (.A0(\register[2] [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27558), .COUT(n27559), .S0(n100[9]), .S1(n100[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_11.INIT0 = 16'h5aaa;
    defparam add_134_11.INIT1 = 16'h5aaa;
    defparam add_134_11.INJECT1_0 = "NO";
    defparam add_134_11.INJECT1_1 = "NO";
    CCU2D add_134_9 (.A0(\register[2] [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27557), .COUT(n27558), .S0(n100[7]), .S1(n100[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_9.INIT0 = 16'h5aaa;
    defparam add_134_9.INIT1 = 16'h5aaa;
    defparam add_134_9.INJECT1_0 = "NO";
    defparam add_134_9.INJECT1_1 = "NO";
    CCU2D add_134_7 (.A0(\register[2] [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27556), .COUT(n27557), .S0(n100[5]), .S1(n100[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_7.INIT0 = 16'h5aaa;
    defparam add_134_7.INIT1 = 16'h5aaa;
    defparam add_134_7.INJECT1_0 = "NO";
    defparam add_134_7.INJECT1_1 = "NO";
    CCU2D add_134_5 (.A0(\register[2][3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27555), .COUT(n27556), .S0(n100[3]), .S1(n100[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_5.INIT0 = 16'h5aaa;
    defparam add_134_5.INIT1 = 16'h5aaa;
    defparam add_134_5.INJECT1_0 = "NO";
    defparam add_134_5.INJECT1_1 = "NO";
    CCU2D add_134_3 (.A0(\register[2] [1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\register[2] [2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27554), .COUT(n27555), .S0(n100[1]), .S1(n100[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_3.INIT0 = 16'h5aaa;
    defparam add_134_3.INIT1 = 16'h5aaa;
    defparam add_134_3.INJECT1_0 = "NO";
    defparam add_134_3.INJECT1_1 = "NO";
    CCU2D add_134_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\register[2][0] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27554), .S1(n100[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(103[23:39])
    defparam add_134_1.INIT0 = 16'hF000;
    defparam add_134_1.INIT1 = 16'h5555;
    defparam add_134_1.INJECT1_0 = "NO";
    defparam add_134_1.INJECT1_1 = "NO";
    \ClockDividerP(factor=12000000)  uptime_div (.debug_c_c(debug_c_c), .clk_1Hz(clk_1Hz), 
            .n32433(n32433), .n34320(n34320), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(107[28] 109[53])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12000000) 
//

module \ClockDividerP(factor=12000000)  (debug_c_c, clk_1Hz, n32433, n34320, 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    output clk_1Hz;
    input n32433;
    input n34320;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n2595;
    wire [31:0]n134;
    
    wire n6778, n30919, n27, n28150, n25, n26, n24, n19, n32, 
        n28, n20, n29, n26_adj_375, n27923, n27922, n27921, n27920, 
        n27919, n27918, n27917, n27916, n27915, n27914, n27913, 
        n27912, n27829, n27828, n27827, n27826, n27825, n27824, 
        n27823, n27822, n27821, n27820, n27819, n27818, n27817, 
        n27816, n27815, n27814;
    
    FD1S3IX count_2175__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2595), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i0.GSR = "ENABLED";
    FD1S3IX clk_o_14 (.D(n6778), .CK(debug_c_c), .CD(n32433), .Q(clk_1Hz));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2175__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2595), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i1.GSR = "ENABLED";
    FD1S3IX count_2175__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2595), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i2.GSR = "ENABLED";
    FD1S3IX count_2175__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2595), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i3.GSR = "ENABLED";
    FD1S3IX count_2175__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2595), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i4.GSR = "ENABLED";
    FD1S3IX count_2175__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2595), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i5.GSR = "ENABLED";
    FD1S3IX count_2175__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2595), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i6.GSR = "ENABLED";
    FD1S3IX count_2175__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2595), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i7.GSR = "ENABLED";
    FD1S3IX count_2175__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2595), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i8.GSR = "ENABLED";
    FD1S3IX count_2175__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2595), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i9.GSR = "ENABLED";
    FD1S3IX count_2175__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i10.GSR = "ENABLED";
    FD1S3IX count_2175__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i11.GSR = "ENABLED";
    FD1S3IX count_2175__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i12.GSR = "ENABLED";
    FD1S3IX count_2175__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i13.GSR = "ENABLED";
    FD1S3IX count_2175__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i14.GSR = "ENABLED";
    FD1S3IX count_2175__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i15.GSR = "ENABLED";
    FD1S3IX count_2175__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i16.GSR = "ENABLED";
    FD1S3IX count_2175__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i17.GSR = "ENABLED";
    FD1S3IX count_2175__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i18.GSR = "ENABLED";
    FD1S3IX count_2175__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i19.GSR = "ENABLED";
    FD1S3IX count_2175__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i20.GSR = "ENABLED";
    FD1S3IX count_2175__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i21.GSR = "ENABLED";
    FD1S3IX count_2175__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i22.GSR = "ENABLED";
    FD1S3IX count_2175__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i23.GSR = "ENABLED";
    FD1S3IX count_2175__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i24.GSR = "ENABLED";
    FD1S3IX count_2175__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i25.GSR = "ENABLED";
    FD1S3IX count_2175__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i26.GSR = "ENABLED";
    FD1S3IX count_2175__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i27.GSR = "ENABLED";
    FD1S3IX count_2175__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i28.GSR = "ENABLED";
    FD1S3IX count_2175__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i29.GSR = "ENABLED";
    FD1S3IX count_2175__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i30.GSR = "ENABLED";
    FD1S3IX count_2175__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2595), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175__i31.GSR = "ENABLED";
    LUT4 i24653_2_lut (.A(n30919), .B(n34320), .Z(n2595)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24653_2_lut.init = 16'heeee;
    LUT4 i24651_4_lut (.A(n27), .B(n28150), .C(n25), .D(n26), .Z(n30919)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i24651_4_lut.init = 16'h0004;
    LUT4 i12_4_lut (.A(count[19]), .B(n24), .C(count[8]), .D(count[14]), 
         .Z(n27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(n19), .B(n32), .C(n28), .D(n20), .Z(n28150)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16_4_lut.init = 16'h8000;
    LUT4 i10_4_lut (.A(count[30]), .B(count[22]), .C(count[13]), .D(count[25]), 
         .Z(n25)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i11_4_lut (.A(count[28]), .B(count[15]), .C(count[31]), .D(count[29]), 
         .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut (.A(count[26]), .B(count[24]), .C(count[10]), .D(count[27]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(29[9:26])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(count[18]), .B(count[1]), .Z(n19)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i15_4_lut (.A(n29), .B(count[9]), .C(n26_adj_375), .D(count[0]), 
         .Z(n32)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i15_4_lut.init = 16'h8000;
    LUT4 i11_4_lut_adj_434 (.A(count[3]), .B(count[12]), .C(count[5]), 
         .D(count[17]), .Z(n28)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i11_4_lut_adj_434.init = 16'h8000;
    LUT4 i3_2_lut (.A(count[2]), .B(count[11]), .Z(n20)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_435 (.A(count[20]), .B(count[7]), .C(count[23]), 
         .D(count[21]), .Z(n29)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12_4_lut_adj_435.init = 16'h8000;
    LUT4 i9_3_lut (.A(count[16]), .B(count[4]), .C(count[6]), .Z(n26_adj_375)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i9_3_lut.init = 16'h8080;
    CCU2D add_21585_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27923), 
          .S0(n6778));
    defparam add_21585_cout.INIT0 = 16'h0000;
    defparam add_21585_cout.INIT1 = 16'h0000;
    defparam add_21585_cout.INJECT1_0 = "NO";
    defparam add_21585_cout.INJECT1_1 = "NO";
    CCU2D add_21585_24 (.A0(count[30]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[31]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27922), .COUT(n27923));
    defparam add_21585_24.INIT0 = 16'h5555;
    defparam add_21585_24.INIT1 = 16'h5555;
    defparam add_21585_24.INJECT1_0 = "NO";
    defparam add_21585_24.INJECT1_1 = "NO";
    CCU2D add_21585_22 (.A0(count[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[29]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27921), .COUT(n27922));
    defparam add_21585_22.INIT0 = 16'h5555;
    defparam add_21585_22.INIT1 = 16'h5555;
    defparam add_21585_22.INJECT1_0 = "NO";
    defparam add_21585_22.INJECT1_1 = "NO";
    CCU2D add_21585_20 (.A0(count[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27920), .COUT(n27921));
    defparam add_21585_20.INIT0 = 16'h5555;
    defparam add_21585_20.INIT1 = 16'h5555;
    defparam add_21585_20.INJECT1_0 = "NO";
    defparam add_21585_20.INJECT1_1 = "NO";
    CCU2D add_21585_18 (.A0(count[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27919), .COUT(n27920));
    defparam add_21585_18.INIT0 = 16'h5555;
    defparam add_21585_18.INIT1 = 16'h5555;
    defparam add_21585_18.INJECT1_0 = "NO";
    defparam add_21585_18.INJECT1_1 = "NO";
    CCU2D add_21585_16 (.A0(count[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27918), .COUT(n27919));
    defparam add_21585_16.INIT0 = 16'h5aaa;
    defparam add_21585_16.INIT1 = 16'h5555;
    defparam add_21585_16.INJECT1_0 = "NO";
    defparam add_21585_16.INJECT1_1 = "NO";
    CCU2D add_21585_14 (.A0(count[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27917), .COUT(n27918));
    defparam add_21585_14.INIT0 = 16'h5aaa;
    defparam add_21585_14.INIT1 = 16'h5555;
    defparam add_21585_14.INJECT1_0 = "NO";
    defparam add_21585_14.INJECT1_1 = "NO";
    CCU2D add_21585_12 (.A0(count[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27916), .COUT(n27917));
    defparam add_21585_12.INIT0 = 16'h5555;
    defparam add_21585_12.INIT1 = 16'h5aaa;
    defparam add_21585_12.INJECT1_0 = "NO";
    defparam add_21585_12.INJECT1_1 = "NO";
    CCU2D add_21585_10 (.A0(count[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27915), .COUT(n27916));
    defparam add_21585_10.INIT0 = 16'h5aaa;
    defparam add_21585_10.INIT1 = 16'h5aaa;
    defparam add_21585_10.INJECT1_0 = "NO";
    defparam add_21585_10.INJECT1_1 = "NO";
    CCU2D add_21585_8 (.A0(count[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27914), .COUT(n27915));
    defparam add_21585_8.INIT0 = 16'h5555;
    defparam add_21585_8.INIT1 = 16'h5aaa;
    defparam add_21585_8.INJECT1_0 = "NO";
    defparam add_21585_8.INJECT1_1 = "NO";
    CCU2D add_21585_6 (.A0(count[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27913), .COUT(n27914));
    defparam add_21585_6.INIT0 = 16'h5555;
    defparam add_21585_6.INIT1 = 16'h5555;
    defparam add_21585_6.INJECT1_0 = "NO";
    defparam add_21585_6.INJECT1_1 = "NO";
    CCU2D add_21585_4 (.A0(count[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27912), .COUT(n27913));
    defparam add_21585_4.INIT0 = 16'h5aaa;
    defparam add_21585_4.INIT1 = 16'h5aaa;
    defparam add_21585_4.INJECT1_0 = "NO";
    defparam add_21585_4.INJECT1_1 = "NO";
    CCU2D add_21585_2 (.A0(count[8]), .B0(count[7]), .C0(GND_net), .D0(GND_net), 
          .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27912));
    defparam add_21585_2.INIT0 = 16'h7000;
    defparam add_21585_2.INIT1 = 16'h5555;
    defparam add_21585_2.INJECT1_0 = "NO";
    defparam add_21585_2.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27829), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_33.INIT1 = 16'h0000;
    defparam count_2175_add_4_33.INJECT1_0 = "NO";
    defparam count_2175_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27828), .COUT(n27829), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_31.INJECT1_0 = "NO";
    defparam count_2175_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27827), .COUT(n27828), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_29.INJECT1_0 = "NO";
    defparam count_2175_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27826), .COUT(n27827), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_27.INJECT1_0 = "NO";
    defparam count_2175_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27825), .COUT(n27826), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_25.INJECT1_0 = "NO";
    defparam count_2175_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27824), .COUT(n27825), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_23.INJECT1_0 = "NO";
    defparam count_2175_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27823), .COUT(n27824), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_21.INJECT1_0 = "NO";
    defparam count_2175_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27822), .COUT(n27823), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_19.INJECT1_0 = "NO";
    defparam count_2175_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27821), .COUT(n27822), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_17.INJECT1_0 = "NO";
    defparam count_2175_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27820), .COUT(n27821), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_15.INJECT1_0 = "NO";
    defparam count_2175_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27819), .COUT(n27820), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_13.INJECT1_0 = "NO";
    defparam count_2175_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27818), .COUT(n27819), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_11.INJECT1_0 = "NO";
    defparam count_2175_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27817), .COUT(n27818), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_9.INJECT1_0 = "NO";
    defparam count_2175_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27816), .COUT(n27817), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_7.INJECT1_0 = "NO";
    defparam count_2175_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27815), .COUT(n27816), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_5.INJECT1_0 = "NO";
    defparam count_2175_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27814), .COUT(n27815), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2175_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2175_add_4_3.INJECT1_0 = "NO";
    defparam count_2175_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2175_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27814), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2175_add_4_1.INIT0 = 16'hF000;
    defparam count_2175_add_4_1.INIT1 = 16'h0555;
    defparam count_2175_add_4_1.INJECT1_0 = "NO";
    defparam count_2175_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0100000) 
//

module \ArmPeripheral(axis_haddr=8'b0100000)  (read_value, debug_c_c, n11981, 
            n32366, \register_addr[1] , n30338, \register_addr[0] , 
            Stepper_Z_M0_c_0, stepping, VCC_net, GND_net, Stepper_Z_nFault_c, 
            n34322, \read_size[0] , n30631, n579, prev_select, n32417, 
            n32505, n32412, n32390, rw, n34320, n32360, databus, 
            n7852, n34323, n608, n610, \control_reg[7] , Stepper_Z_En_c, 
            n34324, Stepper_Z_Dir_c, Stepper_Z_M2_c_2, Stepper_Z_M1_c_1, 
            \read_size[2] , n29663, \steps_reg[5] , \steps_reg[3] , 
            n34325, n28296, n14, n15, n34317, \register_addr[5] , 
            n30310, limit_c_2, \register_addr[4] , n32442, n32503, 
            n32358, n20505, Stepper_Z_Step_c, n32433) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    input n11981;
    input n32366;
    input \register_addr[1] ;
    input n30338;
    input \register_addr[0] ;
    output Stepper_Z_M0_c_0;
    input stepping;
    input VCC_net;
    input GND_net;
    input Stepper_Z_nFault_c;
    input n34322;
    output \read_size[0] ;
    input n30631;
    input n579;
    output prev_select;
    input n32417;
    output n32505;
    input n32412;
    input n32390;
    input rw;
    input n34320;
    input n32360;
    input [31:0]databus;
    input n7852;
    input n34323;
    input n608;
    input n610;
    output \control_reg[7] ;
    output Stepper_Z_En_c;
    input n34324;
    output Stepper_Z_Dir_c;
    output Stepper_Z_M2_c_2;
    output Stepper_Z_M1_c_1;
    output \read_size[2] ;
    input n29663;
    output \steps_reg[5] ;
    output \steps_reg[3] ;
    input n34325;
    output n28296;
    input n14;
    input n15;
    input n34317;
    input \register_addr[5] ;
    input n30310;
    input limit_c_2;
    input \register_addr[4] ;
    input n32442;
    input n32503;
    input n32358;
    output n20505;
    output Stepper_Z_Step_c;
    input n32433;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n30862, n30860, n30861;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire n30339, fault_latched;
    wire [31:0]n3277;
    
    wire n12372, prev_step_clk, step_clk, limit_latched, n182, prev_limit_latched, 
        n12358, n32347, n30818, n30819, n30820;
    wire [31:0]n224;
    
    wire n3276, n9610;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [7:0]n7333;
    wire [31:0]n5746;
    wire [31:0]n5782;
    
    wire n30817, n18847, n6, n30343, n30341, n49, n62, n58, 
        n50, n30344, n30345, n30346, n30347, n30348, n30349, n30350, 
        n30351, n30352, n30342, n30353, n30354, n30355, n30356, 
        n30357, n30358, n30359, n30360, n30361, n30362, n30340, 
        int_step, n20499, n32363, n30815, n30816, n18845, n18848, 
        n5, n27725, n27724, n27723, n27722, n27721, n27720, n27719, 
        n27718, n27717, n27716, n27715, n27714, n27713, n27712, 
        n27711, n27710, n41, n60, n54, n42, n52, n38, n56, 
        n46;
    
    FD1P3IX read_value__i0 (.D(n30862), .SP(n11981), .CD(n32366), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    PFUMX i24503 (.BLUT(n30860), .ALUT(n30861), .C0(\register_addr[1] ), 
          .Z(n30862));
    LUT4 i1_4_lut (.A(div_factor_reg[30]), .B(n30338), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n30339)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i24501_3_lut (.A(Stepper_Z_M0_c_0), .B(stepping), .C(\register_addr[0] ), 
         .Z(n30860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24501_3_lut.init = 16'hcaca;
    IFS1P3DX fault_latched_178 (.D(Stepper_Z_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3277[0]), .CK(debug_c_c), .CD(n34322), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n30631), .SP(n11981), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n12372), .CK(debug_c_c), .Q(Stepper_Z_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n12358), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n32417), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    LUT4 i24502_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n30861)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24502_3_lut.init = 16'hcaca;
    LUT4 i24720_3_lut_rep_253_4_lut_4_lut (.A(n32505), .B(n32412), .C(n32390), 
         .D(rw), .Z(n32347)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i24720_3_lut_rep_253_4_lut_4_lut.init = 16'h0010;
    LUT4 i24742_2_lut_4_lut_4_lut (.A(n32505), .B(n34320), .C(n32360), 
         .D(n32412), .Z(n12372)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i24742_2_lut_4_lut_4_lut.init = 16'hccdc;
    PFUMX i24461 (.BLUT(n30818), .ALUT(n30819), .C0(\register_addr[1] ), 
          .Z(n30820));
    LUT4 mux_1338_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3276), 
         .Z(n3277[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i26_3_lut.init = 16'hcaca;
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n7852), .PD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n7852), .PD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n7852), .PD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n7852), .PD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n7852), .PD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n7852), .PD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n7852), .PD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n12358), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n12358), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n32347), .CD(n9610), .CK(debug_c_c), 
            .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n32347), .PD(n34324), 
            .CK(debug_c_c), .Q(Stepper_Z_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n32347), .PD(n34324), 
            .CK(debug_c_c), .Q(Stepper_Z_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n12372), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n32347), .PD(n34324), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n12372), .CK(debug_c_c), .Q(Stepper_Z_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n32347), .PD(n34324), 
            .CK(debug_c_c), .Q(Stepper_Z_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n29663), .SP(n11981), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    LUT4 mux_1338_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3276), 
         .Z(n3277[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i25_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i31 (.D(n3277[31]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3277[30]), .CK(debug_c_c), .CD(n34322), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3277[29]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3277[28]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3277[27]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3277[26]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3277[25]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3277[24]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3277[23]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3277[22]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3277[21]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3277[20]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3277[19]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3277[18]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3277[17]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3277[16]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3277[15]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3277[14]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3277[13]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3277[12]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3277[11]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3277[10]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3277[9]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3277[8]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3277[7]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3277[6]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3277[5]), .CK(debug_c_c), .CD(n34324), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3277[4]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3277[3]), .CK(debug_c_c), .CD(n34325), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3277[2]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3277[1]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 mux_1338_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3276), 
         .Z(n3277[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3276), 
         .Z(n3277[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3276), 
         .Z(n3277[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3276), 
         .Z(n3277[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3276), 
         .Z(n3277[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3276), 
         .Z(n3277[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3276), 
         .Z(n3277[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3276), 
         .Z(n3277[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3276), 
         .Z(n3277[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3276), 
         .Z(n3277[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3276), 
         .Z(n3277[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3276), 
         .Z(n3277[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3276), 
         .Z(n3277[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i12_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i1 (.D(n30820), .SP(n11981), .CD(n32366), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 mux_1338_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3276), 
         .Z(n3277[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i11_3_lut.init = 16'hcaca;
    LUT4 i13984_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n7333[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13984_2_lut.init = 16'h2222;
    LUT4 mux_1646_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n5746[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1646_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3276), .Z(n3277[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3276), .Z(n3277[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i9_3_lut.init = 16'hcaca;
    PFUMX mux_1650_i5 (.BLUT(n7333[4]), .ALUT(n5746[4]), .C0(\register_addr[1] ), 
          .Z(n5782[4]));
    PFUMX mux_1650_i8 (.BLUT(n7333[7]), .ALUT(n5746[7]), .C0(\register_addr[1] ), 
          .Z(n5782[7]));
    LUT4 mux_1338_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3276), .Z(n3277[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3276), .Z(n3277[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3276), .Z(n3277[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3276), .Z(n3277[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3276), .Z(n3277[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3276), .Z(n3277[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3276), .Z(n3277[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i2_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i2 (.D(n30817), .SP(n11981), .CD(n32366), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n5782[3]), .SP(n11981), .CD(n32366), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n5782[4]), .SP(n11981), .CD(n32366), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n18847), .SP(n11981), .CD(n32366), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6), .SP(n11981), .CD(n32366), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    LUT4 i13982_2_lut (.A(\control_reg[7] ), .B(\register_addr[0] ), .Z(n7333[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13982_2_lut.init = 16'h2222;
    LUT4 mux_1646_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n5746[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1646_i8_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i7 (.D(n5782[7]), .SP(n11981), .CD(n32366), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n30343), .SP(n11981), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n30341), .SP(n11981), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n28296)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    FD1P3AX read_value__i10 (.D(n30344), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n30345), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n30346), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n30347), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n30348), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n30349), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n30350), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n30351), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n30352), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n30342), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n30353), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n30354), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n30355), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n30356), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n30357), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    LUT4 i17_4_lut (.A(steps_reg[0]), .B(steps_reg[9]), .C(steps_reg[28]), 
         .D(steps_reg[2]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    FD1P3AX read_value__i25 (.D(n30358), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n30359), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n30360), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n30361), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n30362), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n30339), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n30340), .SP(n11981), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX int_step_182 (.D(n32363), .SP(n20499), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_411 (.A(div_factor_reg[8]), .B(n30338), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n30343)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_411.init = 16'hc088;
    LUT4 i1_4_lut_adj_412 (.A(div_factor_reg[9]), .B(n30338), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n30341)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_412.init = 16'hc088;
    LUT4 i1_4_lut_adj_413 (.A(div_factor_reg[10]), .B(n30338), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n30344)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_413.init = 16'hc088;
    LUT4 i1_4_lut_adj_414 (.A(div_factor_reg[11]), .B(n30338), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n30345)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_414.init = 16'hc088;
    LUT4 i1_4_lut_adj_415 (.A(div_factor_reg[12]), .B(n30338), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n30346)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_415.init = 16'hc088;
    LUT4 i1_4_lut_adj_416 (.A(div_factor_reg[13]), .B(n30338), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n30347)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_416.init = 16'hc088;
    LUT4 i1_4_lut_adj_417 (.A(div_factor_reg[14]), .B(n30338), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n30348)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_417.init = 16'hc088;
    LUT4 i1_4_lut_adj_418 (.A(div_factor_reg[15]), .B(n30338), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n30349)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_418.init = 16'hc088;
    LUT4 i24456_3_lut (.A(Stepper_Z_M2_c_2), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n30815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24456_3_lut.init = 16'hcaca;
    LUT4 i24457_3_lut (.A(div_factor_reg[2]), .B(steps_reg[2]), .C(\register_addr[0] ), 
         .Z(n30816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24457_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_419 (.A(div_factor_reg[16]), .B(n30338), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n30350)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_419.init = 16'hc088;
    LUT4 i1_4_lut_adj_420 (.A(div_factor_reg[17]), .B(n30338), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n30351)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_420.init = 16'hc088;
    PFUMX i13105 (.BLUT(n18845), .ALUT(n14), .C0(\register_addr[0] ), 
          .Z(n18847));
    PFUMX i13108 (.BLUT(n18848), .ALUT(n15), .C0(\register_addr[0] ), 
          .Z(n5782[3]));
    LUT4 i1_4_lut_adj_421 (.A(div_factor_reg[18]), .B(n30338), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n30352)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_421.init = 16'hc088;
    LUT4 i1_4_lut_adj_422 (.A(div_factor_reg[19]), .B(n30338), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n30342)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_422.init = 16'hc088;
    PFUMX i6 (.BLUT(n7333[6]), .ALUT(n5), .C0(\register_addr[1] ), .Z(n6));
    LUT4 i1_4_lut_adj_423 (.A(div_factor_reg[20]), .B(n30338), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n30353)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_423.init = 16'hc088;
    LUT4 i1_4_lut_adj_424 (.A(div_factor_reg[21]), .B(n30338), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n30354)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_424.init = 16'hc088;
    LUT4 i1_4_lut_adj_425 (.A(div_factor_reg[22]), .B(n30338), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n30355)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_425.init = 16'hc088;
    LUT4 i1_4_lut_adj_426 (.A(div_factor_reg[23]), .B(n30338), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n30356)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_426.init = 16'hc088;
    LUT4 i1_4_lut_adj_427 (.A(div_factor_reg[24]), .B(n30338), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n30357)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_427.init = 16'hc088;
    LUT4 i1_4_lut_adj_428 (.A(div_factor_reg[25]), .B(n30338), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n30358)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_428.init = 16'hc088;
    LUT4 i1_4_lut_adj_429 (.A(div_factor_reg[26]), .B(n30338), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n30359)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_429.init = 16'hc088;
    LUT4 i1_4_lut_adj_430 (.A(div_factor_reg[27]), .B(n30338), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n30360)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_430.init = 16'hc088;
    LUT4 i1_4_lut_adj_431 (.A(div_factor_reg[31]), .B(n30338), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n30340)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_431.init = 16'hc088;
    LUT4 mux_1338_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3276), .Z(n3277[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_432 (.A(div_factor_reg[29]), .B(n30338), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n30362)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_432.init = 16'hc088;
    LUT4 i1_4_lut_adj_433 (.A(div_factor_reg[28]), .B(n30338), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n30361)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_433.init = 16'hc088;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27725), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27724), .COUT(n27725), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27723), .COUT(n27724), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27722), .COUT(n27723), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27721), .COUT(n27722), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27720), .COUT(n27721), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27719), .COUT(n27720), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27718), .COUT(n27719), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27717), .COUT(n27718), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    LUT4 i24459_3_lut (.A(Stepper_Z_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n30818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24459_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27716), .COUT(n27717), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    LUT4 i24460_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n30819)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24460_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27715), .COUT(n27716), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27714), .COUT(n27715), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27713), .COUT(n27714), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27712), .COUT(n27713), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27711), .COUT(n27712), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27710), .COUT(n27711), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(stepping), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n27710), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i3849_3_lut (.A(prev_limit_latched), .B(n34320), .C(limit_latched), 
         .Z(n9610)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i3849_3_lut.init = 16'hdcdc;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_4_lut (.A(n34317), .B(n32390), .C(\register_addr[5] ), 
         .D(n30310), .Z(n3276)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i2_3_lut_4_lut.init = 16'h4000;
    LUT4 i2_3_lut_rep_269 (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .Z(n32363)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i2_3_lut_rep_269.init = 16'h0808;
    LUT4 i14760_4_lut_4_lut (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .D(n34320), .Z(n20499)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i14760_4_lut_4_lut.init = 16'h0038;
    LUT4 i26_4_lut (.A(steps_reg[25]), .B(n52), .C(n38), .D(steps_reg[26]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i118_1_lut (.A(limit_c_2), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i1_2_lut (.A(n7852), .B(n34320), .Z(n12358)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 mux_1338_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3276), 
         .Z(n3277[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i32_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_411 (.A(\register_addr[4] ), .B(\register_addr[5] ), 
         .Z(n32505)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i1_2_lut_rep_411.init = 16'hbbbb;
    LUT4 i18_4_lut (.A(steps_reg[8]), .B(steps_reg[11]), .C(steps_reg[16]), 
         .D(steps_reg[21]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[30]), .B(steps_reg[7]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[20]), .B(n56), .C(n46), .D(steps_reg[15]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[22]), .B(steps_reg[12]), .C(steps_reg[6]), 
         .D(steps_reg[18]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[14]), .B(steps_reg[19]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[13]), .B(steps_reg[17]), .C(\steps_reg[5] ), 
         .D(steps_reg[31]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i13103_3_lut (.A(Stepper_Z_Dir_c), .B(div_factor_reg[5]), .C(\register_addr[1] ), 
         .Z(n18845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13103_3_lut.init = 16'hcaca;
    LUT4 i13106_3_lut (.A(control_reg[3]), .B(div_factor_reg[3]), .C(\register_addr[1] ), 
         .Z(n18848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13106_3_lut.init = 16'hcaca;
    LUT4 i13983_2_lut (.A(Stepper_Z_En_c), .B(\register_addr[0] ), .Z(n7333[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13983_2_lut.init = 16'h2222;
    LUT4 i5_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i5_3_lut.init = 16'hcaca;
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n12358), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=589, LSE_RLINE=602 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 mux_1338_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3276), 
         .Z(n3277[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3276), 
         .Z(n3277[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i30_3_lut.init = 16'hcaca;
    LUT4 i14_2_lut (.A(steps_reg[23]), .B(steps_reg[29]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 mux_1338_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3276), 
         .Z(n3277[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i29_3_lut.init = 16'hcaca;
    LUT4 i24759_2_lut_3_lut_3_lut_4_lut (.A(n32442), .B(n32503), .C(n32358), 
         .D(n34320), .Z(n20505)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i24759_2_lut_3_lut_3_lut_4_lut.init = 16'hff10;
    LUT4 i20_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[27]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(steps_reg[10]), .B(\steps_reg[3] ), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 mux_1338_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3276), 
         .Z(n3277[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1338_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3276), 
         .Z(n3277[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1338_i27_3_lut.init = 16'hcaca;
    LUT4 i24639_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_Z_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i24639_2_lut.init = 16'h9999;
    PFUMX i24458 (.BLUT(n30815), .ALUT(n30816), .C0(\register_addr[1] ), 
          .Z(n30817));
    ClockDivider step_clk_gen (.debug_c_c(debug_c_c), .div_factor_reg({div_factor_reg}), 
            .n34320(n34320), .step_clk(step_clk), .n32433(n32433), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider
//

module ClockDivider (debug_c_c, div_factor_reg, n34320, step_clk, n32433, 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input [31:0]div_factor_reg;
    input n34320;
    output step_clk;
    input n32433;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n32339, n14407, n7056, n7090, n7021;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n27392;
    wire [31:0]n40;
    
    wire n27393, n27391, n27390, n27389, n27388, n27387, n27386, 
        n27385, n27384, n27383, n27382, n27661, n27381, n27380, 
        n27660, n27659, n27379, n27378, n27658, n27657, n27377, 
        n27376, n27656, n27655, n27375, n27654, n27653, n27374, 
        n27373, n27652, n27651, n27372, n27650, n27649, n27371, 
        n27648, n27370, n27647, n27369, n27368, n27646, n27367, 
        n27366, n27365, n27364, n27363, n27362, n27409, n27408, 
        n27407, n27406, n27405, n27404, n27403, n27402, n27401, 
        n27400, n27399, n27398, n27397, n27396, n27395, n27394, 
        n27781, n27780, n27779, n27778, n27777, n27776, n27775, 
        n27774, n27773, n27772, n27771, n27770, n27769, n27768, 
        n27767, n27766;
    
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    LUT4 i962_2_lut_rep_245 (.A(n7056), .B(n34320), .Z(n32339)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i962_2_lut_rep_245.init = 16'heeee;
    LUT4 i8641_2_lut_3_lut (.A(n7056), .B(n34320), .C(n7090), .Z(n14407)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i8641_2_lut_3_lut.init = 16'he0e0;
    FD1S3IX clk_o_22 (.D(n7021), .CK(debug_c_c), .CD(n32433), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    FD1S3IX count_2178__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i0.GSR = "ENABLED";
    FD1S3IX count_2178__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i1.GSR = "ENABLED";
    FD1S3IX count_2178__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i2.GSR = "ENABLED";
    FD1S3IX count_2178__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i3.GSR = "ENABLED";
    FD1S3IX count_2178__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i4.GSR = "ENABLED";
    FD1S3IX count_2178__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i5.GSR = "ENABLED";
    FD1S3IX count_2178__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i6.GSR = "ENABLED";
    FD1S3IX count_2178__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i7.GSR = "ENABLED";
    FD1S3IX count_2178__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i8.GSR = "ENABLED";
    FD1S3IX count_2178__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i9.GSR = "ENABLED";
    FD1S3IX count_2178__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i10.GSR = "ENABLED";
    FD1S3IX count_2178__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i11.GSR = "ENABLED";
    FD1S3IX count_2178__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i12.GSR = "ENABLED";
    FD1S3IX count_2178__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i13.GSR = "ENABLED";
    FD1S3IX count_2178__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i14.GSR = "ENABLED";
    FD1S3IX count_2178__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i15.GSR = "ENABLED";
    FD1S3IX count_2178__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i16.GSR = "ENABLED";
    FD1S3IX count_2178__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i17.GSR = "ENABLED";
    FD1S3IX count_2178__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i18.GSR = "ENABLED";
    FD1S3IX count_2178__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i19.GSR = "ENABLED";
    FD1S3IX count_2178__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i20.GSR = "ENABLED";
    FD1S3IX count_2178__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i21.GSR = "ENABLED";
    FD1S3IX count_2178__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i22.GSR = "ENABLED";
    FD1S3IX count_2178__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i23.GSR = "ENABLED";
    FD1S3IX count_2178__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i24.GSR = "ENABLED";
    FD1S3IX count_2178__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i25.GSR = "ENABLED";
    FD1S3IX count_2178__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i26.GSR = "ENABLED";
    FD1S3IX count_2178__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i27.GSR = "ENABLED";
    FD1S3IX count_2178__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i28.GSR = "ENABLED";
    FD1S3IX count_2178__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i29.GSR = "ENABLED";
    FD1S3IX count_2178__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i30.GSR = "ENABLED";
    FD1S3IX count_2178__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n32339), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178__i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    CCU2D sub_1726_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27392), .COUT(n27393));
    defparam sub_1726_add_2_31.INIT0 = 16'h5999;
    defparam sub_1726_add_2_31.INIT1 = 16'h5999;
    defparam sub_1726_add_2_31.INJECT1_0 = "NO";
    defparam sub_1726_add_2_31.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    CCU2D sub_1726_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27391), .COUT(n27392));
    defparam sub_1726_add_2_29.INIT0 = 16'h5999;
    defparam sub_1726_add_2_29.INIT1 = 16'h5999;
    defparam sub_1726_add_2_29.INJECT1_0 = "NO";
    defparam sub_1726_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27390), .COUT(n27391));
    defparam sub_1726_add_2_27.INIT0 = 16'h5999;
    defparam sub_1726_add_2_27.INIT1 = 16'h5999;
    defparam sub_1726_add_2_27.INJECT1_0 = "NO";
    defparam sub_1726_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27389), .COUT(n27390));
    defparam sub_1726_add_2_25.INIT0 = 16'h5999;
    defparam sub_1726_add_2_25.INIT1 = 16'h5999;
    defparam sub_1726_add_2_25.INJECT1_0 = "NO";
    defparam sub_1726_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27388), .COUT(n27389));
    defparam sub_1726_add_2_23.INIT0 = 16'h5999;
    defparam sub_1726_add_2_23.INIT1 = 16'h5999;
    defparam sub_1726_add_2_23.INJECT1_0 = "NO";
    defparam sub_1726_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27387), .COUT(n27388));
    defparam sub_1726_add_2_21.INIT0 = 16'h5999;
    defparam sub_1726_add_2_21.INIT1 = 16'h5999;
    defparam sub_1726_add_2_21.INJECT1_0 = "NO";
    defparam sub_1726_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27386), .COUT(n27387));
    defparam sub_1726_add_2_19.INIT0 = 16'h5999;
    defparam sub_1726_add_2_19.INIT1 = 16'h5999;
    defparam sub_1726_add_2_19.INJECT1_0 = "NO";
    defparam sub_1726_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27385), .COUT(n27386));
    defparam sub_1726_add_2_17.INIT0 = 16'h5999;
    defparam sub_1726_add_2_17.INIT1 = 16'h5999;
    defparam sub_1726_add_2_17.INJECT1_0 = "NO";
    defparam sub_1726_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27384), .COUT(n27385));
    defparam sub_1726_add_2_15.INIT0 = 16'h5999;
    defparam sub_1726_add_2_15.INIT1 = 16'h5999;
    defparam sub_1726_add_2_15.INJECT1_0 = "NO";
    defparam sub_1726_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27383), .COUT(n27384));
    defparam sub_1726_add_2_13.INIT0 = 16'h5999;
    defparam sub_1726_add_2_13.INIT1 = 16'h5999;
    defparam sub_1726_add_2_13.INJECT1_0 = "NO";
    defparam sub_1726_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27382), .COUT(n27383));
    defparam sub_1726_add_2_11.INIT0 = 16'h5999;
    defparam sub_1726_add_2_11.INIT1 = 16'h5999;
    defparam sub_1726_add_2_11.INJECT1_0 = "NO";
    defparam sub_1726_add_2_11.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27661), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27381), .COUT(n27382));
    defparam sub_1726_add_2_9.INIT0 = 16'h5999;
    defparam sub_1726_add_2_9.INIT1 = 16'h5999;
    defparam sub_1726_add_2_9.INJECT1_0 = "NO";
    defparam sub_1726_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27380), .COUT(n27381));
    defparam sub_1726_add_2_7.INIT0 = 16'h5999;
    defparam sub_1726_add_2_7.INIT1 = 16'h5999;
    defparam sub_1726_add_2_7.INJECT1_0 = "NO";
    defparam sub_1726_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27660), .COUT(n27661), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27659), .COUT(n27660), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27379), .COUT(n27380));
    defparam sub_1726_add_2_5.INIT0 = 16'h5999;
    defparam sub_1726_add_2_5.INIT1 = 16'h5999;
    defparam sub_1726_add_2_5.INJECT1_0 = "NO";
    defparam sub_1726_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27378), .COUT(n27379));
    defparam sub_1726_add_2_3.INIT0 = 16'h5999;
    defparam sub_1726_add_2_3.INIT1 = 16'h5999;
    defparam sub_1726_add_2_3.INJECT1_0 = "NO";
    defparam sub_1726_add_2_3.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27658), .COUT(n27659), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27378));
    defparam sub_1726_add_2_1.INIT0 = 16'h0000;
    defparam sub_1726_add_2_1.INIT1 = 16'h5999;
    defparam sub_1726_add_2_1.INJECT1_0 = "NO";
    defparam sub_1726_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27657), .COUT(n27658), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27377), .S1(n7090));
    defparam sub_1727_add_2_33.INIT0 = 16'hf555;
    defparam sub_1727_add_2_33.INIT1 = 16'h0000;
    defparam sub_1727_add_2_33.INJECT1_0 = "NO";
    defparam sub_1727_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27376), .COUT(n27377));
    defparam sub_1727_add_2_31.INIT0 = 16'hf555;
    defparam sub_1727_add_2_31.INIT1 = 16'hf555;
    defparam sub_1727_add_2_31.INJECT1_0 = "NO";
    defparam sub_1727_add_2_31.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n32339), .CD(n14407), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27656), .COUT(n27657), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27655), .COUT(n27656), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27375), .COUT(n27376));
    defparam sub_1727_add_2_29.INIT0 = 16'hf555;
    defparam sub_1727_add_2_29.INIT1 = 16'hf555;
    defparam sub_1727_add_2_29.INJECT1_0 = "NO";
    defparam sub_1727_add_2_29.INJECT1_1 = "NO";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n32339), .PD(n14407), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27654), .COUT(n27655), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27653), .COUT(n27654), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27374), .COUT(n27375));
    defparam sub_1727_add_2_27.INIT0 = 16'hf555;
    defparam sub_1727_add_2_27.INIT1 = 16'hf555;
    defparam sub_1727_add_2_27.INJECT1_0 = "NO";
    defparam sub_1727_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27373), .COUT(n27374));
    defparam sub_1727_add_2_25.INIT0 = 16'hf555;
    defparam sub_1727_add_2_25.INIT1 = 16'hf555;
    defparam sub_1727_add_2_25.INJECT1_0 = "NO";
    defparam sub_1727_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27652), .COUT(n27653), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27651), .COUT(n27652), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27372), .COUT(n27373));
    defparam sub_1727_add_2_23.INIT0 = 16'hf555;
    defparam sub_1727_add_2_23.INIT1 = 16'hf555;
    defparam sub_1727_add_2_23.INJECT1_0 = "NO";
    defparam sub_1727_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27650), .COUT(n27651), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27649), .COUT(n27650), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27371), .COUT(n27372));
    defparam sub_1727_add_2_21.INIT0 = 16'hf555;
    defparam sub_1727_add_2_21.INIT1 = 16'hf555;
    defparam sub_1727_add_2_21.INJECT1_0 = "NO";
    defparam sub_1727_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27648), .COUT(n27649), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27370), .COUT(n27371));
    defparam sub_1727_add_2_19.INIT0 = 16'hf555;
    defparam sub_1727_add_2_19.INIT1 = 16'hf555;
    defparam sub_1727_add_2_19.INJECT1_0 = "NO";
    defparam sub_1727_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27647), .COUT(n27648), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27369), .COUT(n27370));
    defparam sub_1727_add_2_17.INIT0 = 16'hf555;
    defparam sub_1727_add_2_17.INIT1 = 16'hf555;
    defparam sub_1727_add_2_17.INJECT1_0 = "NO";
    defparam sub_1727_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27368), .COUT(n27369));
    defparam sub_1727_add_2_15.INIT0 = 16'hf555;
    defparam sub_1727_add_2_15.INIT1 = 16'hf555;
    defparam sub_1727_add_2_15.INJECT1_0 = "NO";
    defparam sub_1727_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27646), .COUT(n27647), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27367), .COUT(n27368));
    defparam sub_1727_add_2_13.INIT0 = 16'hf555;
    defparam sub_1727_add_2_13.INIT1 = 16'hf555;
    defparam sub_1727_add_2_13.INJECT1_0 = "NO";
    defparam sub_1727_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27646), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27366), .COUT(n27367));
    defparam sub_1727_add_2_11.INIT0 = 16'hf555;
    defparam sub_1727_add_2_11.INIT1 = 16'hf555;
    defparam sub_1727_add_2_11.INJECT1_0 = "NO";
    defparam sub_1727_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27365), .COUT(n27366));
    defparam sub_1727_add_2_9.INIT0 = 16'hf555;
    defparam sub_1727_add_2_9.INIT1 = 16'hf555;
    defparam sub_1727_add_2_9.INJECT1_0 = "NO";
    defparam sub_1727_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27364), .COUT(n27365));
    defparam sub_1727_add_2_7.INIT0 = 16'hf555;
    defparam sub_1727_add_2_7.INIT1 = 16'hf555;
    defparam sub_1727_add_2_7.INJECT1_0 = "NO";
    defparam sub_1727_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27363), .COUT(n27364));
    defparam sub_1727_add_2_5.INIT0 = 16'hf555;
    defparam sub_1727_add_2_5.INIT1 = 16'hf555;
    defparam sub_1727_add_2_5.INJECT1_0 = "NO";
    defparam sub_1727_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27362), .COUT(n27363));
    defparam sub_1727_add_2_3.INIT0 = 16'hf555;
    defparam sub_1727_add_2_3.INIT1 = 16'hf555;
    defparam sub_1727_add_2_3.INJECT1_0 = "NO";
    defparam sub_1727_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1727_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27362));
    defparam sub_1727_add_2_1.INIT0 = 16'h0000;
    defparam sub_1727_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1727_add_2_1.INJECT1_0 = "NO";
    defparam sub_1727_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27409), .S1(n7021));
    defparam sub_1724_add_2_33.INIT0 = 16'h5555;
    defparam sub_1724_add_2_33.INIT1 = 16'h0000;
    defparam sub_1724_add_2_33.INJECT1_0 = "NO";
    defparam sub_1724_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27408), .COUT(n27409));
    defparam sub_1724_add_2_31.INIT0 = 16'h5999;
    defparam sub_1724_add_2_31.INIT1 = 16'h5999;
    defparam sub_1724_add_2_31.INJECT1_0 = "NO";
    defparam sub_1724_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27407), .COUT(n27408));
    defparam sub_1724_add_2_29.INIT0 = 16'h5999;
    defparam sub_1724_add_2_29.INIT1 = 16'h5999;
    defparam sub_1724_add_2_29.INJECT1_0 = "NO";
    defparam sub_1724_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27406), .COUT(n27407));
    defparam sub_1724_add_2_27.INIT0 = 16'h5999;
    defparam sub_1724_add_2_27.INIT1 = 16'h5999;
    defparam sub_1724_add_2_27.INJECT1_0 = "NO";
    defparam sub_1724_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27405), .COUT(n27406));
    defparam sub_1724_add_2_25.INIT0 = 16'h5999;
    defparam sub_1724_add_2_25.INIT1 = 16'h5999;
    defparam sub_1724_add_2_25.INJECT1_0 = "NO";
    defparam sub_1724_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27404), .COUT(n27405));
    defparam sub_1724_add_2_23.INIT0 = 16'h5999;
    defparam sub_1724_add_2_23.INIT1 = 16'h5999;
    defparam sub_1724_add_2_23.INJECT1_0 = "NO";
    defparam sub_1724_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27403), .COUT(n27404));
    defparam sub_1724_add_2_21.INIT0 = 16'h5999;
    defparam sub_1724_add_2_21.INIT1 = 16'h5999;
    defparam sub_1724_add_2_21.INJECT1_0 = "NO";
    defparam sub_1724_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27402), .COUT(n27403));
    defparam sub_1724_add_2_19.INIT0 = 16'h5999;
    defparam sub_1724_add_2_19.INIT1 = 16'h5999;
    defparam sub_1724_add_2_19.INJECT1_0 = "NO";
    defparam sub_1724_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27401), .COUT(n27402));
    defparam sub_1724_add_2_17.INIT0 = 16'h5999;
    defparam sub_1724_add_2_17.INIT1 = 16'h5999;
    defparam sub_1724_add_2_17.INJECT1_0 = "NO";
    defparam sub_1724_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27400), .COUT(n27401));
    defparam sub_1724_add_2_15.INIT0 = 16'h5999;
    defparam sub_1724_add_2_15.INIT1 = 16'h5999;
    defparam sub_1724_add_2_15.INJECT1_0 = "NO";
    defparam sub_1724_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27399), .COUT(n27400));
    defparam sub_1724_add_2_13.INIT0 = 16'h5999;
    defparam sub_1724_add_2_13.INIT1 = 16'h5999;
    defparam sub_1724_add_2_13.INJECT1_0 = "NO";
    defparam sub_1724_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27398), .COUT(n27399));
    defparam sub_1724_add_2_11.INIT0 = 16'h5999;
    defparam sub_1724_add_2_11.INIT1 = 16'h5999;
    defparam sub_1724_add_2_11.INJECT1_0 = "NO";
    defparam sub_1724_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27397), .COUT(n27398));
    defparam sub_1724_add_2_9.INIT0 = 16'h5999;
    defparam sub_1724_add_2_9.INIT1 = 16'h5999;
    defparam sub_1724_add_2_9.INJECT1_0 = "NO";
    defparam sub_1724_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27396), .COUT(n27397));
    defparam sub_1724_add_2_7.INIT0 = 16'h5999;
    defparam sub_1724_add_2_7.INIT1 = 16'h5999;
    defparam sub_1724_add_2_7.INJECT1_0 = "NO";
    defparam sub_1724_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27395), .COUT(n27396));
    defparam sub_1724_add_2_5.INIT0 = 16'h5999;
    defparam sub_1724_add_2_5.INIT1 = 16'h5999;
    defparam sub_1724_add_2_5.INJECT1_0 = "NO";
    defparam sub_1724_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27394), .COUT(n27395));
    defparam sub_1724_add_2_3.INIT0 = 16'h5999;
    defparam sub_1724_add_2_3.INIT1 = 16'h5999;
    defparam sub_1724_add_2_3.INJECT1_0 = "NO";
    defparam sub_1724_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1724_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27394));
    defparam sub_1724_add_2_1.INIT0 = 16'h0000;
    defparam sub_1724_add_2_1.INIT1 = 16'h5999;
    defparam sub_1724_add_2_1.INJECT1_0 = "NO";
    defparam sub_1724_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1726_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27393), .S1(n7056));
    defparam sub_1726_add_2_33.INIT0 = 16'h5999;
    defparam sub_1726_add_2_33.INIT1 = 16'h0000;
    defparam sub_1726_add_2_33.INJECT1_0 = "NO";
    defparam sub_1726_add_2_33.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27781), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_33.INIT1 = 16'h0000;
    defparam count_2178_add_4_33.INJECT1_0 = "NO";
    defparam count_2178_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27780), .COUT(n27781), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_31.INJECT1_0 = "NO";
    defparam count_2178_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27779), .COUT(n27780), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_29.INJECT1_0 = "NO";
    defparam count_2178_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27778), .COUT(n27779), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_27.INJECT1_0 = "NO";
    defparam count_2178_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27777), .COUT(n27778), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_25.INJECT1_0 = "NO";
    defparam count_2178_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27776), .COUT(n27777), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_23.INJECT1_0 = "NO";
    defparam count_2178_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27775), .COUT(n27776), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_21.INJECT1_0 = "NO";
    defparam count_2178_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27774), .COUT(n27775), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_19.INJECT1_0 = "NO";
    defparam count_2178_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27773), .COUT(n27774), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_17.INJECT1_0 = "NO";
    defparam count_2178_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27772), .COUT(n27773), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_15.INJECT1_0 = "NO";
    defparam count_2178_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27771), .COUT(n27772), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_13.INJECT1_0 = "NO";
    defparam count_2178_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27770), .COUT(n27771), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_11.INJECT1_0 = "NO";
    defparam count_2178_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27769), .COUT(n27770), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_9.INJECT1_0 = "NO";
    defparam count_2178_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27768), .COUT(n27769), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_7.INJECT1_0 = "NO";
    defparam count_2178_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27767), .COUT(n27768), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_5.INJECT1_0 = "NO";
    defparam count_2178_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27766), .COUT(n27767), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2178_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2178_add_4_3.INJECT1_0 = "NO";
    defparam count_2178_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2178_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27766), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2178_add_4_1.INIT0 = 16'hF000;
    defparam count_2178_add_4_1.INIT1 = 16'h0555;
    defparam count_2178_add_4_1.INJECT1_0 = "NO";
    defparam count_2178_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0110000) 
//

module \ArmPeripheral(axis_haddr=8'b0110000)  (read_value, debug_c_c, n12620, 
            GND_net, n30868, register_addr, n32504, n32503, n30240, 
            \steps_reg[0] , n34323, n3181, VCC_net, Stepper_A_nFault_c, 
            \read_size[0] , n30283, Stepper_A_M0_c_0, n20505, n579, 
            div_factor_reg, n12224, prev_select, n32408, n32345, n34321, 
            \databus[31] , \databus[28] , n34322, \databus[13] , \databus[11] , 
            \databus[10] , \databus[9] , \databus[7] , \databus[6] , 
            \databus[5] , n610, \control_reg[7] , Stepper_A_En_c, Stepper_A_Dir_c, 
            \control_reg[4] , \databus[4] , \databus[3] , Stepper_A_M2_c_2, 
            Stepper_A_M1_c_1, \databus[1] , \read_size[2] , n30284, 
            n34324, n34325, \steps_reg[16] , \steps_reg[8] , \steps_reg[5] , 
            \steps_reg[4] , \steps_reg[3] , n32360, n7852, \register[0][2] , 
            force_pause, n21, n32480, n32481, n32440, n32412, n6124, 
            n30211, n17, n224, stepping, n34320, n32454, \register[2][0] , 
            n15, \register[2][3] , n4, n32460, n32442, \div_factor_reg[4] , 
            \div_factor_reg[8] , \databus[8] , \databus[12] , \databus[14] , 
            \databus[15] , \div_factor_reg[16] , \databus[16] , \databus[17] , 
            \databus[18] , \databus[19] , \databus[20] , \databus[21] , 
            \databus[22] , \databus[23] , \databus[24] , \databus[25] , 
            \databus[26] , \databus[27] , \databus[29] , \databus[30] , 
            limit_c_3, Stepper_A_Step_c, n15_adj_187, n28270, n14, 
            n32381, n30427, rw, n32433) /* synthesis syn_module_defined=1 */ ;
    output [31:0]read_value;
    input debug_c_c;
    input n12620;
    input GND_net;
    input n30868;
    input [7:0]register_addr;
    output n32504;
    input n32503;
    output n30240;
    output \steps_reg[0] ;
    input n34323;
    input [31:0]n3181;
    input VCC_net;
    input Stepper_A_nFault_c;
    output \read_size[0] ;
    input n30283;
    output Stepper_A_M0_c_0;
    input n20505;
    input n579;
    output [31:0]div_factor_reg;
    input n12224;
    output prev_select;
    input n32408;
    input n32345;
    input n34321;
    input \databus[31] ;
    input \databus[28] ;
    input n34322;
    input \databus[13] ;
    input \databus[11] ;
    input \databus[10] ;
    input \databus[9] ;
    input \databus[7] ;
    input \databus[6] ;
    input \databus[5] ;
    input n610;
    output \control_reg[7] ;
    output Stepper_A_En_c;
    output Stepper_A_Dir_c;
    output \control_reg[4] ;
    input \databus[4] ;
    input \databus[3] ;
    output Stepper_A_M2_c_2;
    output Stepper_A_M1_c_1;
    input \databus[1] ;
    output \read_size[2] ;
    input n30284;
    input n34324;
    input n34325;
    output \steps_reg[16] ;
    output \steps_reg[8] ;
    output \steps_reg[5] ;
    output \steps_reg[4] ;
    output \steps_reg[3] ;
    input n32360;
    output n7852;
    input \register[0][2] ;
    input force_pause;
    output n21;
    input n32480;
    input n32481;
    output n32440;
    output n32412;
    input n6124;
    input n30211;
    input n17;
    output [31:0]n224;
    input stepping;
    input n34320;
    output n32454;
    input \register[2][0] ;
    output n15;
    input \register[2][3] ;
    output n4;
    output n32460;
    output n32442;
    output \div_factor_reg[4] ;
    output \div_factor_reg[8] ;
    input \databus[8] ;
    input \databus[12] ;
    input \databus[14] ;
    input \databus[15] ;
    output \div_factor_reg[16] ;
    input \databus[16] ;
    input \databus[17] ;
    input \databus[18] ;
    input \databus[19] ;
    input \databus[20] ;
    input \databus[21] ;
    input \databus[22] ;
    input \databus[23] ;
    input \databus[24] ;
    input \databus[25] ;
    input \databus[26] ;
    input \databus[27] ;
    input \databus[29] ;
    input \databus[30] ;
    input limit_c_3;
    output Stepper_A_Step_c;
    input n15_adj_187;
    output n28270;
    input n14;
    input n32381;
    input n30427;
    input rw;
    input n32433;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire n42, fault_latched, prev_step_clk, step_clk, limit_latched, 
        n182, prev_limit_latched;
    wire [31:0]div_factor_reg_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n32346, n9608;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    wire [7:0]n7342;
    wire [31:0]n6060;
    wire [31:0]n6096;
    
    wire n5, n6, n30812, n30813, int_step, n20513, n32361, n30814, 
        n30898, n18809, n30230, n30217, n30218, n30214, n30896, 
        n30897, n18810;
    wire [31:0]n100;
    
    wire n30213, n30215, n30212, n30219, n30220, n30221, n30222, 
        n30223, n30224, n18807, n30225, n30226, n30227, n30228, 
        n30229, n30216, n56, n46, n27709, n27708, n27707, n27706, 
        n27705, n27704, n27703, n27702, n27701, n52, n27700, n27699, 
        n27698, n27697, n27696, n27695, n27694, n38, n49, n62_adj_373, 
        n58, n50, n41, n60_adj_374, n54;
    
    LUT4 i10_2_lut (.A(steps_reg[14]), .B(steps_reg[19]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    FD1P3IX read_value__i0 (.D(n30868), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(register_addr[5]), .B(register_addr[4]), .C(n32504), 
         .D(n32503), .Z(n30240)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i2_4_lut.init = 16'h0002;
    FD1S3IX steps_reg__i0 (.D(n3181[0]), .CK(debug_c_c), .CD(n34323), 
            .Q(\steps_reg[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_A_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n30283), .SP(n12620), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n20505), .CK(debug_c_c), .Q(Stepper_A_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n12224), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n32408), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(\databus[31] ), .SP(n32345), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(\databus[28] ), .SP(n32345), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(\databus[13] ), .SP(n32345), .PD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg_c[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(\databus[11] ), .SP(n32345), .PD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(\databus[10] ), .SP(n32345), .PD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(\databus[9] ), .SP(n32345), .PD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg_c[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(\databus[7] ), .SP(n32345), .PD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg_c[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(\databus[6] ), .SP(n32345), .PD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg_c[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(\databus[5] ), .SP(n32345), .PD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg_c[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n12224), .CK(debug_c_c), 
            .Q(div_factor_reg_c[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(\databus[7] ), .SP(n32346), .CD(n9608), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(\databus[6] ), .SP(n32346), .PD(n34323), 
            .CK(debug_c_c), .Q(Stepper_A_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(\databus[5] ), .SP(n32346), .PD(n34323), 
            .CK(debug_c_c), .Q(Stepper_A_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(\databus[4] ), .SP(n32346), .CD(n34323), 
            .CK(debug_c_c), .Q(\control_reg[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(\databus[3] ), .SP(n32346), .PD(n34323), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n20505), .CK(debug_c_c), .Q(Stepper_A_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(\databus[1] ), .SP(n32346), .PD(n34323), 
            .CK(debug_c_c), .Q(Stepper_A_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n30284), .SP(n12620), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3181[31]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3181[30]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3181[29]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3181[28]), .CK(debug_c_c), .CD(n34321), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3181[27]), .CK(debug_c_c), .CD(n34321), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3181[26]), .CK(debug_c_c), .CD(n34321), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3181[25]), .CK(debug_c_c), .CD(n34321), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3181[24]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3181[23]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3181[22]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3181[21]), .CK(debug_c_c), .CD(n34325), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3181[20]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3181[19]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3181[18]), .CK(debug_c_c), .CD(n34325), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3181[17]), .CK(debug_c_c), .CD(n34325), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3181[16]), .CK(debug_c_c), .CD(n34325), 
            .Q(\steps_reg[16] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3181[15]), .CK(debug_c_c), .CD(n34325), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3181[14]), .CK(debug_c_c), .CD(n34325), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3181[13]), .CK(debug_c_c), .CD(n34325), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3181[12]), .CK(debug_c_c), .CD(n34325), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3181[11]), .CK(debug_c_c), .CD(n34325), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3181[10]), .CK(debug_c_c), .CD(n34325), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3181[9]), .CK(debug_c_c), .CD(n34325), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3181[8]), .CK(debug_c_c), .CD(n34325), 
            .Q(\steps_reg[8] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3181[7]), .CK(debug_c_c), .CD(n34325), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3181[6]), .CK(debug_c_c), .CD(n34325), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3181[5]), .CK(debug_c_c), .CD(n34325), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3181[4]), .CK(debug_c_c), .CD(n34325), 
            .Q(\steps_reg[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3181[3]), .CK(debug_c_c), .CD(n34325), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3181[2]), .CK(debug_c_c), .CD(n34325), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3181[1]), .CK(debug_c_c), .CD(n34325), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 i3_4_lut_4_lut (.A(register_addr[1]), .B(register_addr[0]), .C(n32360), 
         .D(n30240), .Z(n7852)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i3_4_lut_4_lut.init = 16'h2000;
    LUT4 i1_3_lut_4_lut_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(\register[0][2] ), .D(force_pause), .Z(n21)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_3_lut_4_lut_3_lut_4_lut.init = 16'h3332;
    LUT4 i1_2_lut_rep_346_3_lut_4_lut (.A(register_addr[1]), .B(n32504), 
         .C(n32480), .D(n32481), .Z(n32440)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(85[9:13])
    defparam i1_2_lut_rep_346_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_318_3_lut_4_lut (.A(register_addr[1]), .B(n32504), 
         .C(n32503), .D(register_addr[0]), .Z(n32412)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/global.v(85[9:13])
    defparam i1_2_lut_rep_318_3_lut_4_lut.init = 16'hfffe;
    PFUMX mux_1676_i8 (.BLUT(n7342[7]), .ALUT(n6060[7]), .C0(register_addr[1]), 
          .Z(n6096[7]));
    PFUMX i6 (.BLUT(n7342[6]), .ALUT(n5), .C0(register_addr[1]), .Z(n6));
    LUT4 i24453_3_lut (.A(Stepper_A_M1_c_1), .B(fault_latched), .C(register_addr[0]), 
         .Z(n30812)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24453_3_lut.init = 16'hcaca;
    LUT4 i24454_3_lut (.A(div_factor_reg_c[1]), .B(steps_reg[1]), .C(register_addr[0]), 
         .Z(n30813)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24454_3_lut.init = 16'hcaca;
    LUT4 i13973_2_lut (.A(\control_reg[7] ), .B(register_addr[0]), .Z(n7342[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13973_2_lut.init = 16'h2222;
    LUT4 mux_1672_i8_3_lut (.A(div_factor_reg_c[7]), .B(steps_reg[7]), .C(register_addr[0]), 
         .Z(n6060[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1672_i8_3_lut.init = 16'hcaca;
    LUT4 i13974_2_lut (.A(Stepper_A_En_c), .B(register_addr[0]), .Z(n7342[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13974_2_lut.init = 16'h2222;
    LUT4 i5_3_lut (.A(div_factor_reg_c[6]), .B(steps_reg[6]), .C(register_addr[0]), 
         .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i5_3_lut.init = 16'hcaca;
    FD1P3AX int_step_182 (.D(n32361), .SP(n20513), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30814), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30898), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n6096[3]), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n6124), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n18809), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n6096[7]), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n30211), .SP(n12620), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n30230), .SP(n12620), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n30217), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n30218), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n30214), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    LUT4 i24537_3_lut (.A(Stepper_A_M2_c_2), .B(limit_latched), .C(register_addr[0]), 
         .Z(n30896)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24537_3_lut.init = 16'hcaca;
    LUT4 i24538_3_lut (.A(div_factor_reg_c[2]), .B(steps_reg[2]), .C(register_addr[0]), 
         .Z(n30897)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24538_3_lut.init = 16'hcaca;
    LUT4 i13067_3_lut (.A(control_reg[3]), .B(div_factor_reg_c[3]), .C(register_addr[1]), 
         .Z(n18810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13067_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i18 (.D(n100[18]), .SP(n12620), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3IX read_value__i17 (.D(n100[17]), .SP(n12620), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3IX read_value__i16 (.D(n17), .SP(n12620), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3IX read_value__i15 (.D(n100[15]), .SP(n12620), .CD(GND_net), 
            .CK(debug_c_c), .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n30213), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n30215), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n30212), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n30219), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n30220), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n30221), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n30222), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n30223), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n30224), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    LUT4 i13064_3_lut (.A(Stepper_A_Dir_c), .B(div_factor_reg_c[5]), .C(register_addr[1]), 
         .Z(n18807)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13064_3_lut.init = 16'hcaca;
    FD1P3AX read_value__i26 (.D(n30225), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n30226), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n30227), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n30228), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n30229), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n30216), .SP(n12620), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    LUT4 i24_4_lut (.A(steps_reg[13]), .B(steps_reg[17]), .C(\steps_reg[5] ), 
         .D(steps_reg[31]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[23]), .B(steps_reg[29]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i1_4_lut (.A(div_factor_reg_c[9]), .B(register_addr[1]), .C(steps_reg[9]), 
         .D(register_addr[0]), .Z(n30230)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27709), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27708), .COUT(n27709), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27707), .COUT(n27708), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27706), .COUT(n27707), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27705), .COUT(n27706), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27704), .COUT(n27705), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27703), .COUT(n27704), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_392 (.A(div_factor_reg_c[10]), .B(register_addr[1]), 
         .C(steps_reg[10]), .D(register_addr[0]), .Z(n30217)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_392.init = 16'hc088;
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27702), .COUT(n27703), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[16] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27701), .COUT(n27702), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    LUT4 i20_4_lut (.A(steps_reg[24]), .B(\steps_reg[8] ), .C(steps_reg[1]), 
         .D(steps_reg[27]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_393 (.A(div_factor_reg_c[11]), .B(register_addr[1]), 
         .C(steps_reg[11]), .D(register_addr[0]), .Z(n30218)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_393.init = 16'hc088;
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27700), .COUT(n27701), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_394 (.A(div_factor_reg_c[12]), .B(register_addr[1]), 
         .C(steps_reg[12]), .D(register_addr[0]), .Z(n30214)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_394.init = 16'hc088;
    LUT4 i13970_4_lut (.A(div_factor_reg_c[18]), .B(register_addr[1]), .C(steps_reg[18]), 
         .D(register_addr[0]), .Z(n100[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13970_4_lut.init = 16'hc088;
    LUT4 i13971_4_lut (.A(div_factor_reg_c[17]), .B(register_addr[1]), .C(steps_reg[17]), 
         .D(register_addr[0]), .Z(n100[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13971_4_lut.init = 16'hc088;
    LUT4 i2_3_lut_rep_267 (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .Z(n32361)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i2_3_lut_rep_267.init = 16'h0808;
    LUT4 i14774_4_lut_4_lut (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .D(n34320), .Z(n20513)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i14774_4_lut_4_lut.init = 16'h0038;
    LUT4 i13972_4_lut (.A(div_factor_reg_c[15]), .B(register_addr[1]), .C(steps_reg[15]), 
         .D(register_addr[0]), .Z(n100[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13972_4_lut.init = 16'hc088;
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27699), .COUT(n27700), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27698), .COUT(n27699), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[8] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27697), .COUT(n27698), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27696), .COUT(n27697), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\steps_reg[4] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27695), .COUT(n27696), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_395 (.A(div_factor_reg_c[13]), .B(register_addr[1]), 
         .C(steps_reg[13]), .D(register_addr[0]), .Z(n30213)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_395.init = 16'hc088;
    LUT4 i1_4_lut_adj_396 (.A(div_factor_reg_c[14]), .B(register_addr[1]), 
         .C(steps_reg[14]), .D(register_addr[0]), .Z(n30215)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_396.init = 16'hc088;
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27694), .COUT(n27695), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_397 (.A(div_factor_reg_c[19]), .B(register_addr[1]), 
         .C(steps_reg[19]), .D(register_addr[0]), .Z(n30212)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_397.init = 16'hc088;
    LUT4 i1_4_lut_adj_398 (.A(div_factor_reg_c[20]), .B(register_addr[1]), 
         .C(steps_reg[20]), .D(register_addr[0]), .Z(n30219)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_398.init = 16'hc088;
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\steps_reg[0] ), .B1(stepping), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n27694), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_399 (.A(div_factor_reg_c[21]), .B(register_addr[1]), 
         .C(steps_reg[21]), .D(register_addr[0]), .Z(n30220)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_399.init = 16'hc088;
    LUT4 equal_1407_i11_2_lut_rep_410 (.A(register_addr[2]), .B(register_addr[3]), 
         .Z(n32504)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam equal_1407_i11_2_lut_rep_410.init = 16'heeee;
    LUT4 i1_4_lut_adj_400 (.A(div_factor_reg_c[22]), .B(register_addr[1]), 
         .C(steps_reg[22]), .D(register_addr[0]), .Z(n30221)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_400.init = 16'hc088;
    LUT4 i14555_2_lut_rep_360_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[6]), .D(register_addr[7]), .Z(n32454)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i14555_2_lut_rep_360_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut (.A(register_addr[2]), .B(register_addr[3]), .C(\register[2][0] ), 
         .Z(n15)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_4_lut_adj_401 (.A(div_factor_reg_c[23]), .B(register_addr[1]), 
         .C(steps_reg[23]), .D(register_addr[0]), .Z(n30222)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_401.init = 16'hc088;
    LUT4 i1_4_lut_adj_402 (.A(div_factor_reg_c[24]), .B(register_addr[1]), 
         .C(steps_reg[24]), .D(register_addr[0]), .Z(n30223)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_402.init = 16'hc088;
    LUT4 i1_4_lut_adj_403 (.A(div_factor_reg_c[25]), .B(register_addr[1]), 
         .C(steps_reg[25]), .D(register_addr[0]), .Z(n30224)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_403.init = 16'hc088;
    LUT4 i1_2_lut_3_lut_adj_404 (.A(register_addr[2]), .B(register_addr[3]), 
         .C(\register[2][3] ), .Z(n4)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_3_lut_adj_404.init = 16'h1010;
    LUT4 i1_2_lut_rep_366_3_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[1]), .Z(n32460)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_rep_366_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_348_3_lut_4_lut (.A(register_addr[2]), .B(register_addr[3]), 
         .C(register_addr[0]), .D(register_addr[1]), .Z(n32442)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_rep_348_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_405 (.A(div_factor_reg_c[26]), .B(register_addr[1]), 
         .C(steps_reg[26]), .D(register_addr[0]), .Z(n30225)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_405.init = 16'hc088;
    LUT4 i1_4_lut_adj_406 (.A(div_factor_reg_c[27]), .B(register_addr[1]), 
         .C(steps_reg[27]), .D(register_addr[0]), .Z(n30226)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_406.init = 16'hc088;
    LUT4 i6_2_lut (.A(steps_reg[10]), .B(\steps_reg[3] ), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    FD1P3IX div_factor_reg_i1 (.D(\databus[1] ), .SP(n12224), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg_c[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(\databus[3] ), .SP(n12224), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg_c[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(\databus[4] ), .SP(n12224), .CD(n34322), 
            .CK(debug_c_c), .Q(\div_factor_reg[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(\databus[8] ), .SP(n12224), .CD(n34322), 
            .CK(debug_c_c), .Q(\div_factor_reg[8] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(\databus[12] ), .SP(n12224), .CD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg_c[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(\databus[14] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(\databus[15] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(\databus[16] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(\div_factor_reg[16] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(\databus[17] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(\databus[18] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(\databus[19] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(\databus[20] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(\databus[21] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(\databus[22] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(\databus[23] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(\databus[24] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(\databus[25] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(\databus[26] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(\databus[27] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(\databus[29] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(\databus[30] ), .SP(n12224), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg_c[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=604, LSE_RLINE=617 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_407 (.A(div_factor_reg_c[28]), .B(register_addr[1]), 
         .C(steps_reg[28]), .D(register_addr[0]), .Z(n30227)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_407.init = 16'hc088;
    LUT4 i1_4_lut_adj_408 (.A(div_factor_reg_c[29]), .B(register_addr[1]), 
         .C(steps_reg[29]), .D(register_addr[0]), .Z(n30228)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_408.init = 16'hc088;
    LUT4 i1_4_lut_adj_409 (.A(div_factor_reg_c[30]), .B(register_addr[1]), 
         .C(steps_reg[30]), .D(register_addr[0]), .Z(n30229)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_409.init = 16'hc088;
    LUT4 i1_4_lut_adj_410 (.A(div_factor_reg_c[31]), .B(register_addr[1]), 
         .C(steps_reg[31]), .D(register_addr[0]), .Z(n30216)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_410.init = 16'hc088;
    LUT4 i118_1_lut (.A(limit_c_3), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    PFUMX i24455 (.BLUT(n30812), .ALUT(n30813), .C0(register_addr[1]), 
          .Z(n30814));
    LUT4 i3847_3_lut (.A(prev_limit_latched), .B(n34320), .C(limit_latched), 
         .Z(n9608)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i3847_3_lut.init = 16'hdcdc;
    LUT4 i24635_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_A_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i24635_2_lut.init = 16'h9999;
    PFUMX i24539 (.BLUT(n30896), .ALUT(n30897), .C0(register_addr[1]), 
          .Z(n30898));
    PFUMX i13069 (.BLUT(n18810), .ALUT(n15_adj_187), .C0(register_addr[0]), 
          .Z(n6096[3]));
    LUT4 i31_4_lut (.A(n49), .B(n62_adj_373), .C(n58), .D(n50), .Z(n28270)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(\steps_reg[0] ), .B(steps_reg[9]), .C(steps_reg[28]), 
         .D(steps_reg[2]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60_adj_374), .C(n54), .D(n42), .Z(n62_adj_373)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    PFUMX i13066 (.BLUT(n18807), .ALUT(n14), .C0(register_addr[0]), .Z(n18809));
    LUT4 i26_4_lut (.A(steps_reg[25]), .B(n52), .C(n38), .D(steps_reg[26]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(\steps_reg[4] ), .B(steps_reg[11]), .C(\steps_reg[16] ), 
         .D(steps_reg[21]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i24698_2_lut_rep_252_4_lut_4_lut (.A(n32412), .B(n32381), .C(n30427), 
         .D(rw), .Z(n32346)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i24698_2_lut_rep_252_4_lut_4_lut.init = 16'h0040;
    LUT4 i9_2_lut (.A(steps_reg[30]), .B(steps_reg[7]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[20]), .B(n56), .C(n46), .D(steps_reg[15]), 
         .Z(n60_adj_374)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[22]), .B(steps_reg[12]), .C(steps_reg[6]), 
         .D(steps_reg[18]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    ClockDivider_U9 step_clk_gen (.GND_net(GND_net), .debug_c_c(debug_c_c), 
            .div_factor_reg({div_factor_reg_c[31:17], \div_factor_reg[16] , 
            div_factor_reg_c[15:9], \div_factor_reg[8] , div_factor_reg_c[7:5], 
            \div_factor_reg[4] , div_factor_reg_c[3:1], div_factor_reg[0]}), 
            .n34320(n34320), .step_clk(step_clk), .n32433(n32433)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U9
//

module ClockDivider_U9 (GND_net, debug_c_c, div_factor_reg, n34320, 
            step_clk, n32433) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input debug_c_c;
    input [31:0]div_factor_reg;
    input n34320;
    output step_clk;
    input n32433;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n27299;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n27300, n27298, n32340, n14422, n7160, n7194, n7125;
    wire [31:0]n134;
    
    wire n27645;
    wire [31:0]n40;
    
    wire n27644, n27643, n27642, n27641, n27640, n27639, n27638, 
        n27637, n27636, n27635, n27634, n27633, n27632, n27631, 
        n27630, n27308, n27309, n27307, n27306, n27305, n27304, 
        n27313, n27312, n27303, n27311, n27302, n27301, n27310, 
        n27605, n27604, n27603, n27602, n27601, n27600, n27599, 
        n27598, n27597, n27596, n27595, n27594, n27593, n27592, 
        n27591, n27590, n27585, n27584, n27583, n27582, n27581, 
        n27580, n27579, n27578, n27577, n27576, n27575, n27574, 
        n27573, n27572, n27571, n27570, n27813, n27812, n27811, 
        n27810, n27809, n27808, n27807, n27806, n27805, n27804, 
        n27803, n27802, n27801, n27800, n27799, n27798;
    
    CCU2D sub_1729_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27299), .COUT(n27300));
    defparam sub_1729_add_2_5.INIT0 = 16'h5999;
    defparam sub_1729_add_2_5.INIT1 = 16'h5999;
    defparam sub_1729_add_2_5.INJECT1_0 = "NO";
    defparam sub_1729_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27298), .COUT(n27299));
    defparam sub_1729_add_2_3.INIT0 = 16'h5999;
    defparam sub_1729_add_2_3.INIT1 = 16'h5999;
    defparam sub_1729_add_2_3.INJECT1_0 = "NO";
    defparam sub_1729_add_2_3.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    LUT4 i966_2_lut_rep_246 (.A(n7160), .B(n34320), .Z(n32340)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i966_2_lut_rep_246.init = 16'heeee;
    LUT4 i8656_2_lut_3_lut (.A(n7160), .B(n34320), .C(n7194), .Z(n14422)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i8656_2_lut_3_lut.init = 16'he0e0;
    FD1S3IX clk_o_22 (.D(n7125), .CK(debug_c_c), .CD(n32433), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    CCU2D sub_1729_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27298));
    defparam sub_1729_add_2_1.INIT0 = 16'h0000;
    defparam sub_1729_add_2_1.INIT1 = 16'h5999;
    defparam sub_1729_add_2_1.INJECT1_0 = "NO";
    defparam sub_1729_add_2_1.INJECT1_1 = "NO";
    FD1S3IX count_2179__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i0.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1S3IX count_2179__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i1.GSR = "ENABLED";
    FD1S3IX count_2179__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i2.GSR = "ENABLED";
    FD1S3IX count_2179__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i3.GSR = "ENABLED";
    FD1S3IX count_2179__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i4.GSR = "ENABLED";
    FD1S3IX count_2179__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i5.GSR = "ENABLED";
    FD1S3IX count_2179__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i6.GSR = "ENABLED";
    FD1S3IX count_2179__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i7.GSR = "ENABLED";
    FD1S3IX count_2179__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i8.GSR = "ENABLED";
    FD1S3IX count_2179__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i9.GSR = "ENABLED";
    FD1S3IX count_2179__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i10.GSR = "ENABLED";
    FD1S3IX count_2179__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i11.GSR = "ENABLED";
    FD1S3IX count_2179__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i12.GSR = "ENABLED";
    FD1S3IX count_2179__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i13.GSR = "ENABLED";
    FD1S3IX count_2179__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i14.GSR = "ENABLED";
    FD1S3IX count_2179__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i15.GSR = "ENABLED";
    FD1S3IX count_2179__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i16.GSR = "ENABLED";
    FD1S3IX count_2179__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i17.GSR = "ENABLED";
    FD1S3IX count_2179__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i18.GSR = "ENABLED";
    FD1S3IX count_2179__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i19.GSR = "ENABLED";
    FD1S3IX count_2179__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i20.GSR = "ENABLED";
    FD1S3IX count_2179__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i21.GSR = "ENABLED";
    FD1S3IX count_2179__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i22.GSR = "ENABLED";
    FD1S3IX count_2179__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i23.GSR = "ENABLED";
    FD1S3IX count_2179__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i24.GSR = "ENABLED";
    FD1S3IX count_2179__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i25.GSR = "ENABLED";
    FD1S3IX count_2179__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i26.GSR = "ENABLED";
    FD1S3IX count_2179__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i27.GSR = "ENABLED";
    FD1S3IX count_2179__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i28.GSR = "ENABLED";
    FD1S3IX count_2179__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i29.GSR = "ENABLED";
    FD1S3IX count_2179__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i30.GSR = "ENABLED";
    FD1S3IX count_2179__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n32340), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179__i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n32340), .CD(n14422), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n32340), .PD(n14422), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27645), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27644), .COUT(n27645), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27643), .COUT(n27644), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27642), .COUT(n27643), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27641), .COUT(n27642), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27640), .COUT(n27641), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27639), .COUT(n27640), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27638), .COUT(n27639), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27637), .COUT(n27638), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27636), .COUT(n27637), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27635), .COUT(n27636), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27634), .COUT(n27635), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27633), .COUT(n27634), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27632), .COUT(n27633), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27631), .COUT(n27632), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27630), .COUT(n27631), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27630), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27308), .COUT(n27309));
    defparam sub_1729_add_2_23.INIT0 = 16'h5999;
    defparam sub_1729_add_2_23.INIT1 = 16'h5999;
    defparam sub_1729_add_2_23.INJECT1_0 = "NO";
    defparam sub_1729_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27307), .COUT(n27308));
    defparam sub_1729_add_2_21.INIT0 = 16'h5999;
    defparam sub_1729_add_2_21.INIT1 = 16'h5999;
    defparam sub_1729_add_2_21.INJECT1_0 = "NO";
    defparam sub_1729_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27306), .COUT(n27307));
    defparam sub_1729_add_2_19.INIT0 = 16'h5999;
    defparam sub_1729_add_2_19.INIT1 = 16'h5999;
    defparam sub_1729_add_2_19.INJECT1_0 = "NO";
    defparam sub_1729_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27305), .COUT(n27306));
    defparam sub_1729_add_2_17.INIT0 = 16'h5999;
    defparam sub_1729_add_2_17.INIT1 = 16'h5999;
    defparam sub_1729_add_2_17.INJECT1_0 = "NO";
    defparam sub_1729_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27304), .COUT(n27305));
    defparam sub_1729_add_2_15.INIT0 = 16'h5999;
    defparam sub_1729_add_2_15.INIT1 = 16'h5999;
    defparam sub_1729_add_2_15.INJECT1_0 = "NO";
    defparam sub_1729_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27313), .S1(n7125));
    defparam sub_1729_add_2_33.INIT0 = 16'h5555;
    defparam sub_1729_add_2_33.INIT1 = 16'h0000;
    defparam sub_1729_add_2_33.INJECT1_0 = "NO";
    defparam sub_1729_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27312), .COUT(n27313));
    defparam sub_1729_add_2_31.INIT0 = 16'h5999;
    defparam sub_1729_add_2_31.INIT1 = 16'h5999;
    defparam sub_1729_add_2_31.INJECT1_0 = "NO";
    defparam sub_1729_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27303), .COUT(n27304));
    defparam sub_1729_add_2_13.INIT0 = 16'h5999;
    defparam sub_1729_add_2_13.INIT1 = 16'h5999;
    defparam sub_1729_add_2_13.INJECT1_0 = "NO";
    defparam sub_1729_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27311), .COUT(n27312));
    defparam sub_1729_add_2_29.INIT0 = 16'h5999;
    defparam sub_1729_add_2_29.INIT1 = 16'h5999;
    defparam sub_1729_add_2_29.INJECT1_0 = "NO";
    defparam sub_1729_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27302), .COUT(n27303));
    defparam sub_1729_add_2_11.INIT0 = 16'h5999;
    defparam sub_1729_add_2_11.INIT1 = 16'h5999;
    defparam sub_1729_add_2_11.INJECT1_0 = "NO";
    defparam sub_1729_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27301), .COUT(n27302));
    defparam sub_1729_add_2_9.INIT0 = 16'h5999;
    defparam sub_1729_add_2_9.INIT1 = 16'h5999;
    defparam sub_1729_add_2_9.INJECT1_0 = "NO";
    defparam sub_1729_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27310), .COUT(n27311));
    defparam sub_1729_add_2_27.INIT0 = 16'h5999;
    defparam sub_1729_add_2_27.INIT1 = 16'h5999;
    defparam sub_1729_add_2_27.INJECT1_0 = "NO";
    defparam sub_1729_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27300), .COUT(n27301));
    defparam sub_1729_add_2_7.INIT0 = 16'h5999;
    defparam sub_1729_add_2_7.INIT1 = 16'h5999;
    defparam sub_1729_add_2_7.INJECT1_0 = "NO";
    defparam sub_1729_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1729_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27309), .COUT(n27310));
    defparam sub_1729_add_2_25.INIT0 = 16'h5999;
    defparam sub_1729_add_2_25.INIT1 = 16'h5999;
    defparam sub_1729_add_2_25.INJECT1_0 = "NO";
    defparam sub_1729_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27605), .S1(n7160));
    defparam sub_1731_add_2_33.INIT0 = 16'h5999;
    defparam sub_1731_add_2_33.INIT1 = 16'h0000;
    defparam sub_1731_add_2_33.INJECT1_0 = "NO";
    defparam sub_1731_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27604), .COUT(n27605));
    defparam sub_1731_add_2_31.INIT0 = 16'h5999;
    defparam sub_1731_add_2_31.INIT1 = 16'h5999;
    defparam sub_1731_add_2_31.INJECT1_0 = "NO";
    defparam sub_1731_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27603), .COUT(n27604));
    defparam sub_1731_add_2_29.INIT0 = 16'h5999;
    defparam sub_1731_add_2_29.INIT1 = 16'h5999;
    defparam sub_1731_add_2_29.INJECT1_0 = "NO";
    defparam sub_1731_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27602), .COUT(n27603));
    defparam sub_1731_add_2_27.INIT0 = 16'h5999;
    defparam sub_1731_add_2_27.INIT1 = 16'h5999;
    defparam sub_1731_add_2_27.INJECT1_0 = "NO";
    defparam sub_1731_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27601), .COUT(n27602));
    defparam sub_1731_add_2_25.INIT0 = 16'h5999;
    defparam sub_1731_add_2_25.INIT1 = 16'h5999;
    defparam sub_1731_add_2_25.INJECT1_0 = "NO";
    defparam sub_1731_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27600), .COUT(n27601));
    defparam sub_1731_add_2_23.INIT0 = 16'h5999;
    defparam sub_1731_add_2_23.INIT1 = 16'h5999;
    defparam sub_1731_add_2_23.INJECT1_0 = "NO";
    defparam sub_1731_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27599), .COUT(n27600));
    defparam sub_1731_add_2_21.INIT0 = 16'h5999;
    defparam sub_1731_add_2_21.INIT1 = 16'h5999;
    defparam sub_1731_add_2_21.INJECT1_0 = "NO";
    defparam sub_1731_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27598), .COUT(n27599));
    defparam sub_1731_add_2_19.INIT0 = 16'h5999;
    defparam sub_1731_add_2_19.INIT1 = 16'h5999;
    defparam sub_1731_add_2_19.INJECT1_0 = "NO";
    defparam sub_1731_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27597), .COUT(n27598));
    defparam sub_1731_add_2_17.INIT0 = 16'h5999;
    defparam sub_1731_add_2_17.INIT1 = 16'h5999;
    defparam sub_1731_add_2_17.INJECT1_0 = "NO";
    defparam sub_1731_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27596), .COUT(n27597));
    defparam sub_1731_add_2_15.INIT0 = 16'h5999;
    defparam sub_1731_add_2_15.INIT1 = 16'h5999;
    defparam sub_1731_add_2_15.INJECT1_0 = "NO";
    defparam sub_1731_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27595), .COUT(n27596));
    defparam sub_1731_add_2_13.INIT0 = 16'h5999;
    defparam sub_1731_add_2_13.INIT1 = 16'h5999;
    defparam sub_1731_add_2_13.INJECT1_0 = "NO";
    defparam sub_1731_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27594), .COUT(n27595));
    defparam sub_1731_add_2_11.INIT0 = 16'h5999;
    defparam sub_1731_add_2_11.INIT1 = 16'h5999;
    defparam sub_1731_add_2_11.INJECT1_0 = "NO";
    defparam sub_1731_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27593), .COUT(n27594));
    defparam sub_1731_add_2_9.INIT0 = 16'h5999;
    defparam sub_1731_add_2_9.INIT1 = 16'h5999;
    defparam sub_1731_add_2_9.INJECT1_0 = "NO";
    defparam sub_1731_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27592), .COUT(n27593));
    defparam sub_1731_add_2_7.INIT0 = 16'h5999;
    defparam sub_1731_add_2_7.INIT1 = 16'h5999;
    defparam sub_1731_add_2_7.INJECT1_0 = "NO";
    defparam sub_1731_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27591), .COUT(n27592));
    defparam sub_1731_add_2_5.INIT0 = 16'h5999;
    defparam sub_1731_add_2_5.INIT1 = 16'h5999;
    defparam sub_1731_add_2_5.INJECT1_0 = "NO";
    defparam sub_1731_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27590), .COUT(n27591));
    defparam sub_1731_add_2_3.INIT0 = 16'h5999;
    defparam sub_1731_add_2_3.INIT1 = 16'h5999;
    defparam sub_1731_add_2_3.INJECT1_0 = "NO";
    defparam sub_1731_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1731_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27590));
    defparam sub_1731_add_2_1.INIT0 = 16'h0000;
    defparam sub_1731_add_2_1.INIT1 = 16'h5999;
    defparam sub_1731_add_2_1.INJECT1_0 = "NO";
    defparam sub_1731_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27585), .S1(n7194));
    defparam sub_1732_add_2_33.INIT0 = 16'hf555;
    defparam sub_1732_add_2_33.INIT1 = 16'h0000;
    defparam sub_1732_add_2_33.INJECT1_0 = "NO";
    defparam sub_1732_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27584), .COUT(n27585));
    defparam sub_1732_add_2_31.INIT0 = 16'hf555;
    defparam sub_1732_add_2_31.INIT1 = 16'hf555;
    defparam sub_1732_add_2_31.INJECT1_0 = "NO";
    defparam sub_1732_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27583), .COUT(n27584));
    defparam sub_1732_add_2_29.INIT0 = 16'hf555;
    defparam sub_1732_add_2_29.INIT1 = 16'hf555;
    defparam sub_1732_add_2_29.INJECT1_0 = "NO";
    defparam sub_1732_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27582), .COUT(n27583));
    defparam sub_1732_add_2_27.INIT0 = 16'hf555;
    defparam sub_1732_add_2_27.INIT1 = 16'hf555;
    defparam sub_1732_add_2_27.INJECT1_0 = "NO";
    defparam sub_1732_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27581), .COUT(n27582));
    defparam sub_1732_add_2_25.INIT0 = 16'hf555;
    defparam sub_1732_add_2_25.INIT1 = 16'hf555;
    defparam sub_1732_add_2_25.INJECT1_0 = "NO";
    defparam sub_1732_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27580), .COUT(n27581));
    defparam sub_1732_add_2_23.INIT0 = 16'hf555;
    defparam sub_1732_add_2_23.INIT1 = 16'hf555;
    defparam sub_1732_add_2_23.INJECT1_0 = "NO";
    defparam sub_1732_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27579), .COUT(n27580));
    defparam sub_1732_add_2_21.INIT0 = 16'hf555;
    defparam sub_1732_add_2_21.INIT1 = 16'hf555;
    defparam sub_1732_add_2_21.INJECT1_0 = "NO";
    defparam sub_1732_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27578), .COUT(n27579));
    defparam sub_1732_add_2_19.INIT0 = 16'hf555;
    defparam sub_1732_add_2_19.INIT1 = 16'hf555;
    defparam sub_1732_add_2_19.INJECT1_0 = "NO";
    defparam sub_1732_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27577), .COUT(n27578));
    defparam sub_1732_add_2_17.INIT0 = 16'hf555;
    defparam sub_1732_add_2_17.INIT1 = 16'hf555;
    defparam sub_1732_add_2_17.INJECT1_0 = "NO";
    defparam sub_1732_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27576), .COUT(n27577));
    defparam sub_1732_add_2_15.INIT0 = 16'hf555;
    defparam sub_1732_add_2_15.INIT1 = 16'hf555;
    defparam sub_1732_add_2_15.INJECT1_0 = "NO";
    defparam sub_1732_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27575), .COUT(n27576));
    defparam sub_1732_add_2_13.INIT0 = 16'hf555;
    defparam sub_1732_add_2_13.INIT1 = 16'hf555;
    defparam sub_1732_add_2_13.INJECT1_0 = "NO";
    defparam sub_1732_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27574), .COUT(n27575));
    defparam sub_1732_add_2_11.INIT0 = 16'hf555;
    defparam sub_1732_add_2_11.INIT1 = 16'hf555;
    defparam sub_1732_add_2_11.INJECT1_0 = "NO";
    defparam sub_1732_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27573), .COUT(n27574));
    defparam sub_1732_add_2_9.INIT0 = 16'hf555;
    defparam sub_1732_add_2_9.INIT1 = 16'hf555;
    defparam sub_1732_add_2_9.INJECT1_0 = "NO";
    defparam sub_1732_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27572), .COUT(n27573));
    defparam sub_1732_add_2_7.INIT0 = 16'hf555;
    defparam sub_1732_add_2_7.INIT1 = 16'hf555;
    defparam sub_1732_add_2_7.INJECT1_0 = "NO";
    defparam sub_1732_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27571), .COUT(n27572));
    defparam sub_1732_add_2_5.INIT0 = 16'hf555;
    defparam sub_1732_add_2_5.INIT1 = 16'hf555;
    defparam sub_1732_add_2_5.INJECT1_0 = "NO";
    defparam sub_1732_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27570), .COUT(n27571));
    defparam sub_1732_add_2_3.INIT0 = 16'hf555;
    defparam sub_1732_add_2_3.INIT1 = 16'hf555;
    defparam sub_1732_add_2_3.INJECT1_0 = "NO";
    defparam sub_1732_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1732_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27570));
    defparam sub_1732_add_2_1.INIT0 = 16'h0000;
    defparam sub_1732_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1732_add_2_1.INJECT1_0 = "NO";
    defparam sub_1732_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27813), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_33.INIT1 = 16'h0000;
    defparam count_2179_add_4_33.INJECT1_0 = "NO";
    defparam count_2179_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27812), .COUT(n27813), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_31.INJECT1_0 = "NO";
    defparam count_2179_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27811), .COUT(n27812), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_29.INJECT1_0 = "NO";
    defparam count_2179_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27810), .COUT(n27811), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_27.INJECT1_0 = "NO";
    defparam count_2179_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27809), .COUT(n27810), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_25.INJECT1_0 = "NO";
    defparam count_2179_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27808), .COUT(n27809), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_23.INJECT1_0 = "NO";
    defparam count_2179_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27807), .COUT(n27808), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_21.INJECT1_0 = "NO";
    defparam count_2179_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27806), .COUT(n27807), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_19.INJECT1_0 = "NO";
    defparam count_2179_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27805), .COUT(n27806), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_17.INJECT1_0 = "NO";
    defparam count_2179_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27804), .COUT(n27805), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_15.INJECT1_0 = "NO";
    defparam count_2179_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27803), .COUT(n27804), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_13.INJECT1_0 = "NO";
    defparam count_2179_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27802), .COUT(n27803), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_11.INJECT1_0 = "NO";
    defparam count_2179_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27801), .COUT(n27802), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_9.INJECT1_0 = "NO";
    defparam count_2179_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27800), .COUT(n27801), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_7.INJECT1_0 = "NO";
    defparam count_2179_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27799), .COUT(n27800), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_5.INJECT1_0 = "NO";
    defparam count_2179_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27798), .COUT(n27799), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2179_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2179_add_4_3.INJECT1_0 = "NO";
    defparam count_2179_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2179_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27798), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2179_add_4_1.INIT0 = 16'hF000;
    defparam count_2179_add_4_1.INIT1 = 16'h0555;
    defparam count_2179_add_4_1.INJECT1_0 = "NO";
    defparam count_2179_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b010000) 
//

module \ArmPeripheral(axis_haddr=8'b010000)  (databus, n3363, debug_c_c, 
            n34322, VCC_net, GND_net, Stepper_Y_nFault_c, \read_size[0] , 
            n30710, Stepper_Y_M0_c_0, n579, \register_addr[5] , \register_addr[4] , 
            n11883, n12434, \arm_select[1] , read_value, n32504, n32503, 
            n32480, \select[4] , n32401, n32348, n34321, n34324, 
            n34323, n34325, \control_reg[7] , Stepper_Y_En_c, Stepper_Y_Dir_c, 
            Stepper_Y_M2_c_2, Stepper_Y_M1_c_1, \read_size[2] , n30411, 
            n30427, n32408, n32505, n32417, n34326, \steps_reg[5] , 
            \steps_reg[3] , limit_c_1, stepping, \register_addr[0] , 
            n34320, \register_addr[1] , n14, n15, n28309, n32412, 
            n32389, rw, Stepper_Y_Step_c, n52, n34317, n32365, n32433) /* synthesis syn_module_defined=1 */ ;
    input [31:0]databus;
    input n3363;
    input debug_c_c;
    input n34322;
    input VCC_net;
    input GND_net;
    input Stepper_Y_nFault_c;
    output \read_size[0] ;
    input n30710;
    output Stepper_Y_M0_c_0;
    input n579;
    input \register_addr[5] ;
    input \register_addr[4] ;
    output n11883;
    input n12434;
    input \arm_select[1] ;
    output [31:0]read_value;
    input n32504;
    input n32503;
    input n32480;
    input \select[4] ;
    output n32401;
    input n32348;
    input n34321;
    input n34324;
    input n34323;
    input n34325;
    output \control_reg[7] ;
    output Stepper_Y_En_c;
    output Stepper_Y_Dir_c;
    output Stepper_Y_M2_c_2;
    output Stepper_Y_M1_c_1;
    output \read_size[2] ;
    input n30411;
    input n30427;
    output n32408;
    input n32505;
    output n32417;
    input n34326;
    output \steps_reg[5] ;
    output \steps_reg[3] ;
    input limit_c_1;
    input stepping;
    input \register_addr[0] ;
    input n34320;
    input \register_addr[1] ;
    input n14;
    input n15;
    output n28309;
    input n32412;
    output n32389;
    input rw;
    output Stepper_Y_Step_c;
    output n52;
    input n34317;
    output n32365;
    input n32433;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]n224;
    wire [31:0]n3364;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire fault_latched, n12954, n20491, prev_step_clk, step_clk, limit_latched, 
        n182, prev_limit_latched;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire prev_select, n30859, n32364, n9612;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n30857, n30858, int_step, n20503, n32359;
    wire [7:0]n7324;
    wire [31:0]n5432;
    
    wire n30821, n30822, n30823, n18883, n18885, n27741, n27740, 
        n18886;
    wire [31:0]n5468;
    
    wire n27739, n27738, n27737, n30824, n30825, n30826, n27736, 
        n27735, n5, n6, n27734, n27733, n27732, n27731, n27730, 
        n27729, n27728, n27727, n49, n62, n58, n50, n27726, 
        n41, n60, n54, n42, n52_c, n38, n56, n46, n32416, 
        n30287, n30294, n30295, n30296, n30297, n30303, n30286, 
        n30293, n30298, n30299, n30288, n30305, n30301, n30308, 
        n30292, n30302, n30290, n30291, n30304, n30289, n30306, 
        n30309, n30300, n30307;
    
    LUT4 mux_1361_i1_3_lut (.A(n224[0]), .B(databus[0]), .C(n3363), .Z(n3364[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i1_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i0 (.D(n3364[0]), .CK(debug_c_c), .CD(n34322), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_Y_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    FD1P3AX read_size__i1 (.D(n30710), .SP(n12954), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n20491), .CK(debug_c_c), .Q(Stepper_Y_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(\register_addr[5] ), .B(\register_addr[4] ), .Z(n11883)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i1_2_lut.init = 16'hbbbb;
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n12434), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(\arm_select[1] ), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1P3IX read_value__i0 (.D(n30859), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_307_3_lut_4_lut (.A(n32504), .B(n32503), .C(n32480), 
         .D(\select[4] ), .Z(n32401)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_307_3_lut_4_lut.init = 16'h0100;
    FD1P3JX div_factor_reg_i13 (.D(databus[13]), .SP(n32348), .PD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(databus[11]), .SP(n32348), .PD(n34324), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(databus[10]), .SP(n32348), .PD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(databus[9]), .SP(n32348), .PD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i8 (.D(databus[8]), .SP(n32348), .CD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(databus[7]), .SP(n32348), .PD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(databus[6]), .SP(n32348), .PD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(databus[5]), .SP(n32348), .PD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i4 (.D(databus[4]), .SP(n32348), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(databus[3]), .SP(n32348), .CD(n34323), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i2 (.D(databus[2]), .SP(n32348), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i1 (.D(databus[1]), .SP(n32348), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(databus[7]), .SP(n32364), .CD(n9612), .CK(debug_c_c), 
            .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(databus[6]), .SP(n32364), .PD(n34325), 
            .CK(debug_c_c), .Q(Stepper_Y_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(databus[5]), .SP(n32364), .PD(n34325), 
            .CK(debug_c_c), .Q(Stepper_Y_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3IX control_reg_i5 (.D(databus[4]), .SP(n32364), .CD(n34321), 
            .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(databus[3]), .SP(n32364), .PD(n34325), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3IX control_reg_i3 (.D(databus[2]), .SP(n32364), .CD(n34325), 
            .CK(debug_c_c), .Q(Stepper_Y_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(databus[1]), .SP(n32364), .PD(n34325), 
            .CK(debug_c_c), .Q(Stepper_Y_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n30411), .SP(n12954), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_314_3_lut_4_lut (.A(n32504), .B(n32503), .C(n30427), 
         .D(\select[4] ), .Z(n32408)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_314_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_323_3_lut_4_lut (.A(n32504), .B(n32503), .C(n32505), 
         .D(\select[4] ), .Z(n32417)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_323_3_lut_4_lut.init = 16'h0100;
    FD1S3IX steps_reg__i31 (.D(n3364[31]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    FD1S3IX steps_reg__i30 (.D(n3364[30]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3364[29]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3364[28]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3364[27]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3364[26]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3364[25]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3364[24]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3364[23]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3364[22]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3364[21]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3364[20]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    FD1S3IX steps_reg__i19 (.D(n3364[19]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    FD1S3IX steps_reg__i18 (.D(n3364[18]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    FD1S3IX steps_reg__i17 (.D(n3364[17]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3364[16]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3364[15]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3364[14]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3364[13]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3364[12]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3364[11]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3364[10]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3364[9]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3364[8]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3364[7]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3364[6]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3364[5]), .CK(debug_c_c), .CD(n34326), 
            .Q(\steps_reg[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3364[4]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3364[3]), .CK(debug_c_c), .CD(n34326), 
            .Q(\steps_reg[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3364[2]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3364[1]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    LUT4 i118_1_lut (.A(limit_c_1), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    LUT4 i24498_3_lut (.A(Stepper_Y_M0_c_0), .B(stepping), .C(\register_addr[0] ), 
         .Z(n30857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24498_3_lut.init = 16'hcaca;
    LUT4 i24499_3_lut (.A(div_factor_reg[0]), .B(steps_reg[0]), .C(\register_addr[0] ), 
         .Z(n30858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24499_3_lut.init = 16'hcaca;
    LUT4 i3851_3_lut (.A(prev_limit_latched), .B(n34320), .C(limit_latched), 
         .Z(n9612)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i3851_3_lut.init = 16'hdcdc;
    LUT4 mux_1361_i32_3_lut (.A(n224[31]), .B(databus[31]), .C(n3363), 
         .Z(n3364[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i32_3_lut.init = 16'hcaca;
    FD1P3AX int_step_182 (.D(n32359), .SP(n20503), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    LUT4 i13987_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n7324[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13987_2_lut.init = 16'h2222;
    LUT4 mux_1620_i5_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n5432[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1620_i5_3_lut.init = 16'hcaca;
    LUT4 i13985_2_lut (.A(\control_reg[7] ), .B(\register_addr[0] ), .Z(n7324[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13985_2_lut.init = 16'h2222;
    LUT4 mux_1620_i8_3_lut (.A(div_factor_reg[7]), .B(steps_reg[7]), .C(\register_addr[0] ), 
         .Z(n5432[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1620_i8_3_lut.init = 16'hcaca;
    PFUMX i24464 (.BLUT(n30821), .ALUT(n30822), .C0(\register_addr[1] ), 
          .Z(n30823));
    PFUMX i13144 (.BLUT(n18883), .ALUT(n14), .C0(\register_addr[0] ), 
          .Z(n18885));
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27741), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27740), .COUT(n27741), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    PFUMX i13147 (.BLUT(n18886), .ALUT(n15), .C0(\register_addr[0] ), 
          .Z(n5468[3]));
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27739), .COUT(n27740), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27738), .COUT(n27739), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27737), .COUT(n27738), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    PFUMX i24467 (.BLUT(n30824), .ALUT(n30825), .C0(\register_addr[1] ), 
          .Z(n30826));
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27736), .COUT(n27737), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27735), .COUT(n27736), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    PFUMX i6 (.BLUT(n7324[6]), .ALUT(n5), .C0(\register_addr[1] ), .Z(n6));
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27734), .COUT(n27735), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27733), .COUT(n27734), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27732), .COUT(n27733), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27731), .COUT(n27732), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27730), .COUT(n27731), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    LUT4 mux_1361_i31_3_lut (.A(n224[30]), .B(databus[30]), .C(n3363), 
         .Z(n3364[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i31_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_9 (.A0(steps_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27729), .COUT(n27730), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    LUT4 mux_1361_i30_3_lut (.A(n224[29]), .B(databus[29]), .C(n3363), 
         .Z(n3364[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i30_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_7 (.A0(\steps_reg[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27728), .COUT(n27729), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    LUT4 mux_1361_i29_3_lut (.A(n224[28]), .B(databus[28]), .C(n3363), 
         .Z(n3364[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i29_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_5 (.A0(\steps_reg[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27727), .COUT(n27728), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    LUT4 mux_1361_i28_3_lut (.A(n224[27]), .B(databus[27]), .C(n3363), 
         .Z(n3364[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i27_3_lut (.A(n224[26]), .B(databus[26]), .C(n3363), 
         .Z(n3364[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i27_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n28309)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 mux_1361_i26_3_lut (.A(n224[25]), .B(databus[25]), .C(n3363), 
         .Z(n3364[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i26_3_lut.init = 16'hcaca;
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27726), .COUT(n27727), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    LUT4 i17_4_lut (.A(steps_reg[0]), .B(steps_reg[9]), .C(steps_reg[28]), 
         .D(steps_reg[2]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 mux_1361_i25_3_lut (.A(n224[24]), .B(databus[24]), .C(n3363), 
         .Z(n3364[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i25_3_lut.init = 16'hcaca;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[25]), .B(n52_c), .C(n38), .D(steps_reg[26]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(stepping), .C1(step_clk), .D1(prev_step_clk), 
          .COUT(n27726), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    LUT4 i18_4_lut (.A(steps_reg[8]), .B(steps_reg[11]), .C(steps_reg[16]), 
         .D(steps_reg[21]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 mux_1361_i24_3_lut (.A(n224[23]), .B(databus[23]), .C(n3363), 
         .Z(n3364[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i23_3_lut (.A(n224[22]), .B(databus[22]), .C(n3363), 
         .Z(n3364[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i22_3_lut (.A(n224[21]), .B(databus[21]), .C(n3363), 
         .Z(n3364[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i22_3_lut.init = 16'hcaca;
    LUT4 i9_2_lut (.A(steps_reg[30]), .B(steps_reg[7]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[20]), .B(n56), .C(n46), .D(steps_reg[15]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(steps_reg[22]), .B(steps_reg[12]), .C(steps_reg[6]), 
         .D(steps_reg[18]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[14]), .B(steps_reg[19]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 mux_1361_i21_3_lut (.A(n224[20]), .B(databus[20]), .C(n3363), 
         .Z(n3364[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i20_3_lut (.A(n224[19]), .B(databus[19]), .C(n3363), 
         .Z(n3364[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i20_3_lut.init = 16'hcaca;
    LUT4 i24_4_lut (.A(steps_reg[13]), .B(steps_reg[17]), .C(\steps_reg[5] ), 
         .D(steps_reg[31]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[23]), .B(steps_reg[29]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 mux_1361_i19_3_lut (.A(n224[18]), .B(databus[18]), .C(n3363), 
         .Z(n3364[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i18_3_lut (.A(n224[17]), .B(databus[17]), .C(n3363), 
         .Z(n3364[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i18_3_lut.init = 16'hcaca;
    LUT4 i20_4_lut (.A(steps_reg[24]), .B(steps_reg[4]), .C(steps_reg[1]), 
         .D(steps_reg[27]), .Z(n52_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 mux_1361_i17_3_lut (.A(n224[16]), .B(databus[16]), .C(n3363), 
         .Z(n3364[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i16_3_lut (.A(n224[15]), .B(databus[15]), .C(n3363), 
         .Z(n3364[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i15_3_lut (.A(n224[14]), .B(databus[14]), .C(n3363), 
         .Z(n3364[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i14_3_lut (.A(n224[13]), .B(databus[13]), .C(n3363), 
         .Z(n3364[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i13_3_lut (.A(n224[12]), .B(databus[12]), .C(n3363), 
         .Z(n3364[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i12_3_lut (.A(n224[11]), .B(databus[11]), .C(n3363), 
         .Z(n3364[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i11_3_lut (.A(n224[10]), .B(databus[10]), .C(n3363), 
         .Z(n3364[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i10_3_lut (.A(n224[9]), .B(databus[9]), .C(n3363), .Z(n3364[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i9_3_lut (.A(n224[8]), .B(databus[8]), .C(n3363), .Z(n3364[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i8_3_lut (.A(n224[7]), .B(databus[7]), .C(n3363), .Z(n3364[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i7_3_lut (.A(n224[6]), .B(databus[6]), .C(n3363), .Z(n3364[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i6_3_lut (.A(n224[5]), .B(databus[5]), .C(n3363), .Z(n3364[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i5_3_lut (.A(n224[4]), .B(databus[4]), .C(n3363), .Z(n3364[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i4_3_lut (.A(n224[3]), .B(databus[3]), .C(n3363), .Z(n3364[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i3_3_lut (.A(n224[2]), .B(databus[2]), .C(n3363), .Z(n3364[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1361_i2_3_lut (.A(n224[1]), .B(databus[1]), .C(n3363), .Z(n3364[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam mux_1361_i2_3_lut.init = 16'hcaca;
    LUT4 i6_2_lut (.A(steps_reg[10]), .B(\steps_reg[3] ), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i24704_2_lut_4_lut_4_lut (.A(n32412), .B(n34320), .C(n11883), 
         .D(n32389), .Z(n20491)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(118[11:28])
    defparam i24704_2_lut_4_lut_4_lut.init = 16'hcdcc;
    LUT4 i2_3_lut_rep_265 (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .Z(n32359)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i2_3_lut_rep_265.init = 16'h0808;
    LUT4 i14764_4_lut_4_lut (.A(stepping), .B(step_clk), .C(prev_step_clk), 
         .D(n34320), .Z(n20503)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(76[9:45])
    defparam i14764_4_lut_4_lut.init = 16'h0038;
    FD1P3IX div_factor_reg_i12 (.D(databus[12]), .SP(n12434), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(databus[14]), .SP(n12434), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i15 (.D(databus[15]), .SP(n12434), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i16 (.D(databus[16]), .SP(n12434), .CD(n34324), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(databus[17]), .SP(n12434), .CD(n34324), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(databus[18]), .SP(n12434), .CD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(databus[19]), .SP(n12434), .CD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(databus[20]), .SP(n12434), .CD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(databus[21]), .SP(n12434), .CD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(databus[22]), .SP(n12434), .CD(n34324), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(databus[23]), .SP(n12434), .CD(n34324), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(databus[24]), .SP(n12434), .CD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(databus[25]), .SP(n12434), .CD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(databus[26]), .SP(n12434), .CD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(databus[27]), .SP(n12434), .CD(n34322), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(databus[28]), .SP(n12434), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(databus[29]), .SP(n12434), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(databus[30]), .SP(n12434), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(databus[31]), .SP(n12434), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    LUT4 i24462_3_lut (.A(Stepper_Y_M2_c_2), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n30821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24462_3_lut.init = 16'hcaca;
    LUT4 i24463_3_lut (.A(div_factor_reg[2]), .B(steps_reg[2]), .C(\register_addr[0] ), 
         .Z(n30822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24463_3_lut.init = 16'hcaca;
    LUT4 i13142_3_lut (.A(Stepper_Y_Dir_c), .B(div_factor_reg[5]), .C(\register_addr[1] ), 
         .Z(n18883)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13142_3_lut.init = 16'hcaca;
    LUT4 i13145_3_lut (.A(control_reg[3]), .B(div_factor_reg[3]), .C(\register_addr[1] ), 
         .Z(n18886)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i13145_3_lut.init = 16'hcaca;
    LUT4 i24465_3_lut (.A(Stepper_Y_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n30824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24465_3_lut.init = 16'hcaca;
    LUT4 i24466_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n30825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24466_3_lut.init = 16'hcaca;
    LUT4 i13986_2_lut (.A(Stepper_Y_En_c), .B(\register_addr[0] ), .Z(n7324[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i13986_2_lut.init = 16'h2222;
    LUT4 i5_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), .C(\register_addr[0] ), 
         .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i5_3_lut.init = 16'hcaca;
    LUT4 i24711_3_lut_rep_270_3_lut_4_lut (.A(rw), .B(n32416), .C(n11883), 
         .D(n32412), .Z(n32364)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i24711_3_lut_rep_270_3_lut_4_lut.init = 16'h0004;
    FD1P3AX read_value__i31 (.D(n30287), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n30294), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n30295), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n30296), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n30297), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n30303), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n30286), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n30293), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n30298), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n30299), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n30288), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n30305), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n30301), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n30308), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n30292), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n30302), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i15 (.D(n30290), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n30291), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n30304), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n30289), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i11 (.D(n30306), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n30309), .SP(n12954), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    FD1P3AX read_value__i9 (.D(n30300), .SP(n12954), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n30307), .SP(n12954), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n5468[7]), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n6), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n18885), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n5468[4]), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX read_value__i3 (.D(n5468[3]), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX read_value__i2 (.D(n30823), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30826), .SP(n12954), .CD(GND_net), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=574, LSE_RLINE=587 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    PFUMX i24500 (.BLUT(n30857), .ALUT(n30858), .C0(\register_addr[1] ), 
          .Z(n30859));
    LUT4 i1_4_lut (.A(div_factor_reg[31]), .B(\register_addr[1] ), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n30287)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_369 (.A(div_factor_reg[30]), .B(\register_addr[1] ), 
         .C(steps_reg[30]), .D(\register_addr[0] ), .Z(n30294)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_369.init = 16'hc088;
    LUT4 i1_4_lut_adj_370 (.A(div_factor_reg[29]), .B(\register_addr[1] ), 
         .C(steps_reg[29]), .D(\register_addr[0] ), .Z(n30295)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_370.init = 16'hc088;
    LUT4 i1_4_lut_adj_371 (.A(div_factor_reg[28]), .B(\register_addr[1] ), 
         .C(steps_reg[28]), .D(\register_addr[0] ), .Z(n30296)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_371.init = 16'hc088;
    LUT4 i24641_2_lut (.A(int_step), .B(control_reg[3]), .Z(Stepper_Y_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    defparam i24641_2_lut.init = 16'h9999;
    LUT4 i20_2_lut (.A(\arm_select[1] ), .B(rw), .Z(n52)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(55[19:32])
    defparam i20_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_372 (.A(div_factor_reg[27]), .B(\register_addr[1] ), 
         .C(steps_reg[27]), .D(\register_addr[0] ), .Z(n30297)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_372.init = 16'hc088;
    LUT4 i1_4_lut_adj_373 (.A(div_factor_reg[26]), .B(\register_addr[1] ), 
         .C(steps_reg[26]), .D(\register_addr[0] ), .Z(n30303)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_373.init = 16'hc088;
    LUT4 i1_4_lut_adj_374 (.A(div_factor_reg[25]), .B(\register_addr[1] ), 
         .C(steps_reg[25]), .D(\register_addr[0] ), .Z(n30286)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_374.init = 16'hc088;
    PFUMX mux_1624_i5 (.BLUT(n7324[4]), .ALUT(n5432[4]), .C0(\register_addr[1] ), 
          .Z(n5468[4]));
    LUT4 i1_4_lut_adj_375 (.A(div_factor_reg[24]), .B(\register_addr[1] ), 
         .C(steps_reg[24]), .D(\register_addr[0] ), .Z(n30293)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_375.init = 16'hc088;
    LUT4 i1_4_lut_adj_376 (.A(div_factor_reg[23]), .B(\register_addr[1] ), 
         .C(steps_reg[23]), .D(\register_addr[0] ), .Z(n30298)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_376.init = 16'hc088;
    PFUMX mux_1624_i8 (.BLUT(n7324[7]), .ALUT(n5432[7]), .C0(\register_addr[1] ), 
          .Z(n5468[7]));
    LUT4 i1_4_lut_adj_377 (.A(div_factor_reg[22]), .B(\register_addr[1] ), 
         .C(steps_reg[22]), .D(\register_addr[0] ), .Z(n30299)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_377.init = 16'hc088;
    LUT4 i1_4_lut_adj_378 (.A(div_factor_reg[21]), .B(\register_addr[1] ), 
         .C(steps_reg[21]), .D(\register_addr[0] ), .Z(n30288)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_378.init = 16'hc088;
    LUT4 i1_4_lut_adj_379 (.A(div_factor_reg[20]), .B(\register_addr[1] ), 
         .C(steps_reg[20]), .D(\register_addr[0] ), .Z(n30305)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_379.init = 16'hc088;
    LUT4 i1_4_lut_adj_380 (.A(div_factor_reg[19]), .B(\register_addr[1] ), 
         .C(steps_reg[19]), .D(\register_addr[0] ), .Z(n30301)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_380.init = 16'hc088;
    LUT4 i1_4_lut_adj_381 (.A(div_factor_reg[18]), .B(\register_addr[1] ), 
         .C(steps_reg[18]), .D(\register_addr[0] ), .Z(n30308)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_381.init = 16'hc088;
    LUT4 i1_4_lut_adj_382 (.A(div_factor_reg[17]), .B(\register_addr[1] ), 
         .C(steps_reg[17]), .D(\register_addr[0] ), .Z(n30292)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_382.init = 16'hc088;
    LUT4 i1_2_lut_rep_322 (.A(\arm_select[1] ), .B(prev_select), .Z(n32416)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i1_2_lut_rep_322.init = 16'h2222;
    LUT4 i1_4_lut_adj_383 (.A(div_factor_reg[16]), .B(\register_addr[1] ), 
         .C(steps_reg[16]), .D(\register_addr[0] ), .Z(n30302)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_383.init = 16'hc088;
    LUT4 i1_4_lut_adj_384 (.A(div_factor_reg[15]), .B(\register_addr[1] ), 
         .C(steps_reg[15]), .D(\register_addr[0] ), .Z(n30290)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_384.init = 16'hc088;
    LUT4 i1_4_lut_adj_385 (.A(div_factor_reg[14]), .B(\register_addr[1] ), 
         .C(steps_reg[14]), .D(\register_addr[0] ), .Z(n30291)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_385.init = 16'hc088;
    LUT4 i1_4_lut_adj_386 (.A(div_factor_reg[13]), .B(\register_addr[1] ), 
         .C(steps_reg[13]), .D(\register_addr[0] ), .Z(n30304)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_386.init = 16'hc088;
    LUT4 i1_2_lut_rep_295_3_lut (.A(\arm_select[1] ), .B(prev_select), .C(n34317), 
         .Z(n32389)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i1_2_lut_rep_295_3_lut.init = 16'h0202;
    LUT4 i1_2_lut_rep_271_3_lut_4_lut (.A(\arm_select[1] ), .B(prev_select), 
         .C(\register_addr[5] ), .D(rw), .Z(n32365)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i1_2_lut_rep_271_3_lut_4_lut.init = 16'h0002;
    LUT4 i1_4_lut_adj_387 (.A(div_factor_reg[12]), .B(\register_addr[1] ), 
         .C(steps_reg[12]), .D(\register_addr[0] ), .Z(n30289)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_387.init = 16'hc088;
    LUT4 i1_2_lut_2_lut_3_lut (.A(\arm_select[1] ), .B(prev_select), .C(n34320), 
         .Z(n12954)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i1_2_lut_2_lut_3_lut.init = 16'h0202;
    LUT4 i1_4_lut_adj_388 (.A(div_factor_reg[11]), .B(\register_addr[1] ), 
         .C(steps_reg[11]), .D(\register_addr[0] ), .Z(n30306)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_388.init = 16'hc088;
    LUT4 i1_4_lut_adj_389 (.A(div_factor_reg[10]), .B(\register_addr[1] ), 
         .C(steps_reg[10]), .D(\register_addr[0] ), .Z(n30309)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_389.init = 16'hc088;
    LUT4 i1_4_lut_adj_390 (.A(div_factor_reg[9]), .B(\register_addr[1] ), 
         .C(steps_reg[9]), .D(\register_addr[0] ), .Z(n30300)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_390.init = 16'hc088;
    LUT4 i1_4_lut_adj_391 (.A(div_factor_reg[8]), .B(\register_addr[1] ), 
         .C(steps_reg[8]), .D(\register_addr[0] ), .Z(n30307)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_391.init = 16'hc088;
    ClockDivider_U7 step_clk_gen (.debug_c_c(debug_c_c), .div_factor_reg({div_factor_reg}), 
            .n34320(n34320), .step_clk(step_clk), .n32433(n32433), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U7
//

module ClockDivider_U7 (debug_c_c, div_factor_reg, n34320, step_clk, 
            n32433, GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input [31:0]div_factor_reg;
    input n34320;
    output step_clk;
    input n32433;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    
    wire n32338, n14396, n6952, n6986, n6917;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n27677;
    wire [31:0]n40;
    
    wire n27676, n27675, n27674, n27673, n27672, n27671, n27670, 
        n27669, n27668, n27667, n27666, n27665, n27664, n27663, 
        n27662, n27457, n27456, n27455, n27454, n27453, n27452, 
        n27451, n27450, n27449, n27448, n27447, n27446, n27445, 
        n27444, n27443, n27442, n27441, n27440, n27439, n27438, 
        n27437, n27436, n27435, n27434, n27433, n27432, n27431, 
        n27430, n27429, n27428, n27427, n27426, n27425, n27424, 
        n27423, n27422, n27421, n27420, n27419, n27418, n27417, 
        n27416, n27415, n27414, n27413, n27412, n27411, n27410, 
        n27877, n27876, n27875, n27874, n27873, n27872, n27871, 
        n27870, n27869, n27868, n27867, n27866, n27865, n27864, 
        n27863, n27862;
    
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    LUT4 i8630_2_lut_3_lut (.A(n6952), .B(n34320), .C(n6986), .Z(n14396)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i8630_2_lut_3_lut.init = 16'he0e0;
    LUT4 i958_2_lut_rep_244 (.A(n6952), .B(n34320), .Z(n32338)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i958_2_lut_rep_244.init = 16'heeee;
    FD1S3IX clk_o_22 (.D(n6917), .CK(debug_c_c), .CD(n32433), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    FD1S3IX count_2177__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i0.GSR = "ENABLED";
    FD1S3IX count_2177__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i1.GSR = "ENABLED";
    FD1S3IX count_2177__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i2.GSR = "ENABLED";
    FD1S3IX count_2177__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i3.GSR = "ENABLED";
    FD1S3IX count_2177__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i4.GSR = "ENABLED";
    FD1S3IX count_2177__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i5.GSR = "ENABLED";
    FD1S3IX count_2177__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i6.GSR = "ENABLED";
    FD1S3IX count_2177__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i7.GSR = "ENABLED";
    FD1S3IX count_2177__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i8.GSR = "ENABLED";
    FD1S3IX count_2177__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i9.GSR = "ENABLED";
    FD1S3IX count_2177__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i10.GSR = "ENABLED";
    FD1S3IX count_2177__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i11.GSR = "ENABLED";
    FD1S3IX count_2177__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i12.GSR = "ENABLED";
    FD1S3IX count_2177__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i13.GSR = "ENABLED";
    FD1S3IX count_2177__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i14.GSR = "ENABLED";
    FD1S3IX count_2177__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i15.GSR = "ENABLED";
    FD1S3IX count_2177__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i16.GSR = "ENABLED";
    FD1S3IX count_2177__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i17.GSR = "ENABLED";
    FD1S3IX count_2177__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i18.GSR = "ENABLED";
    FD1S3IX count_2177__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i19.GSR = "ENABLED";
    FD1S3IX count_2177__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i20.GSR = "ENABLED";
    FD1S3IX count_2177__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i21.GSR = "ENABLED";
    FD1S3IX count_2177__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i22.GSR = "ENABLED";
    FD1S3IX count_2177__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i23.GSR = "ENABLED";
    FD1S3IX count_2177__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i24.GSR = "ENABLED";
    FD1S3IX count_2177__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i25.GSR = "ENABLED";
    FD1S3IX count_2177__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i26.GSR = "ENABLED";
    FD1S3IX count_2177__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i27.GSR = "ENABLED";
    FD1S3IX count_2177__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i28.GSR = "ENABLED";
    FD1S3IX count_2177__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i29.GSR = "ENABLED";
    FD1S3IX count_2177__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i30.GSR = "ENABLED";
    FD1S3IX count_2177__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n32338), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177__i31.GSR = "ENABLED";
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27677), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27676), .COUT(n27677), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27675), .COUT(n27676), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27674), .COUT(n27675), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27673), .COUT(n27674), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27672), .COUT(n27673), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27671), .COUT(n27672), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27670), .COUT(n27671), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27669), .COUT(n27670), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27668), .COUT(n27669), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27667), .COUT(n27668), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27666), .COUT(n27667), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27665), .COUT(n27666), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27664), .COUT(n27665), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27663), .COUT(n27664), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27662), .COUT(n27663), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27662), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    CCU2D sub_1719_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27457), .S1(n6917));
    defparam sub_1719_add_2_33.INIT0 = 16'h5555;
    defparam sub_1719_add_2_33.INIT1 = 16'h0000;
    defparam sub_1719_add_2_33.INJECT1_0 = "NO";
    defparam sub_1719_add_2_33.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    CCU2D sub_1719_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27456), .COUT(n27457));
    defparam sub_1719_add_2_31.INIT0 = 16'h5999;
    defparam sub_1719_add_2_31.INIT1 = 16'h5999;
    defparam sub_1719_add_2_31.INJECT1_0 = "NO";
    defparam sub_1719_add_2_31.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    CCU2D sub_1719_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27455), .COUT(n27456));
    defparam sub_1719_add_2_29.INIT0 = 16'h5999;
    defparam sub_1719_add_2_29.INIT1 = 16'h5999;
    defparam sub_1719_add_2_29.INJECT1_0 = "NO";
    defparam sub_1719_add_2_29.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    CCU2D sub_1719_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27454), .COUT(n27455));
    defparam sub_1719_add_2_27.INIT0 = 16'h5999;
    defparam sub_1719_add_2_27.INIT1 = 16'h5999;
    defparam sub_1719_add_2_27.INJECT1_0 = "NO";
    defparam sub_1719_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27453), .COUT(n27454));
    defparam sub_1719_add_2_25.INIT0 = 16'h5999;
    defparam sub_1719_add_2_25.INIT1 = 16'h5999;
    defparam sub_1719_add_2_25.INJECT1_0 = "NO";
    defparam sub_1719_add_2_25.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    CCU2D sub_1719_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27452), .COUT(n27453));
    defparam sub_1719_add_2_23.INIT0 = 16'h5999;
    defparam sub_1719_add_2_23.INIT1 = 16'h5999;
    defparam sub_1719_add_2_23.INJECT1_0 = "NO";
    defparam sub_1719_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27451), .COUT(n27452));
    defparam sub_1719_add_2_21.INIT0 = 16'h5999;
    defparam sub_1719_add_2_21.INIT1 = 16'h5999;
    defparam sub_1719_add_2_21.INJECT1_0 = "NO";
    defparam sub_1719_add_2_21.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    CCU2D sub_1719_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27450), .COUT(n27451));
    defparam sub_1719_add_2_19.INIT0 = 16'h5999;
    defparam sub_1719_add_2_19.INIT1 = 16'h5999;
    defparam sub_1719_add_2_19.INJECT1_0 = "NO";
    defparam sub_1719_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27449), .COUT(n27450));
    defparam sub_1719_add_2_17.INIT0 = 16'h5999;
    defparam sub_1719_add_2_17.INIT1 = 16'h5999;
    defparam sub_1719_add_2_17.INJECT1_0 = "NO";
    defparam sub_1719_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27448), .COUT(n27449));
    defparam sub_1719_add_2_15.INIT0 = 16'h5999;
    defparam sub_1719_add_2_15.INIT1 = 16'h5999;
    defparam sub_1719_add_2_15.INJECT1_0 = "NO";
    defparam sub_1719_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27447), .COUT(n27448));
    defparam sub_1719_add_2_13.INIT0 = 16'h5999;
    defparam sub_1719_add_2_13.INIT1 = 16'h5999;
    defparam sub_1719_add_2_13.INJECT1_0 = "NO";
    defparam sub_1719_add_2_13.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    CCU2D sub_1719_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27446), .COUT(n27447));
    defparam sub_1719_add_2_11.INIT0 = 16'h5999;
    defparam sub_1719_add_2_11.INIT1 = 16'h5999;
    defparam sub_1719_add_2_11.INJECT1_0 = "NO";
    defparam sub_1719_add_2_11.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    CCU2D sub_1719_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27445), .COUT(n27446));
    defparam sub_1719_add_2_9.INIT0 = 16'h5999;
    defparam sub_1719_add_2_9.INIT1 = 16'h5999;
    defparam sub_1719_add_2_9.INJECT1_0 = "NO";
    defparam sub_1719_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27444), .COUT(n27445));
    defparam sub_1719_add_2_7.INIT0 = 16'h5999;
    defparam sub_1719_add_2_7.INIT1 = 16'h5999;
    defparam sub_1719_add_2_7.INJECT1_0 = "NO";
    defparam sub_1719_add_2_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n32338), .CD(n14396), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    CCU2D sub_1719_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27443), .COUT(n27444));
    defparam sub_1719_add_2_5.INIT0 = 16'h5999;
    defparam sub_1719_add_2_5.INIT1 = 16'h5999;
    defparam sub_1719_add_2_5.INJECT1_0 = "NO";
    defparam sub_1719_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27442), .COUT(n27443));
    defparam sub_1719_add_2_3.INIT0 = 16'h5999;
    defparam sub_1719_add_2_3.INIT1 = 16'h5999;
    defparam sub_1719_add_2_3.INJECT1_0 = "NO";
    defparam sub_1719_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1719_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27442));
    defparam sub_1719_add_2_1.INIT0 = 16'h0000;
    defparam sub_1719_add_2_1.INIT1 = 16'h5999;
    defparam sub_1719_add_2_1.INJECT1_0 = "NO";
    defparam sub_1719_add_2_1.INJECT1_1 = "NO";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n32338), .PD(n14396), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    CCU2D sub_1721_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27441), .S1(n6952));
    defparam sub_1721_add_2_33.INIT0 = 16'h5999;
    defparam sub_1721_add_2_33.INIT1 = 16'h0000;
    defparam sub_1721_add_2_33.INJECT1_0 = "NO";
    defparam sub_1721_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27440), .COUT(n27441));
    defparam sub_1721_add_2_31.INIT0 = 16'h5999;
    defparam sub_1721_add_2_31.INIT1 = 16'h5999;
    defparam sub_1721_add_2_31.INJECT1_0 = "NO";
    defparam sub_1721_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27439), .COUT(n27440));
    defparam sub_1721_add_2_29.INIT0 = 16'h5999;
    defparam sub_1721_add_2_29.INIT1 = 16'h5999;
    defparam sub_1721_add_2_29.INJECT1_0 = "NO";
    defparam sub_1721_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27438), .COUT(n27439));
    defparam sub_1721_add_2_27.INIT0 = 16'h5999;
    defparam sub_1721_add_2_27.INIT1 = 16'h5999;
    defparam sub_1721_add_2_27.INJECT1_0 = "NO";
    defparam sub_1721_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27437), .COUT(n27438));
    defparam sub_1721_add_2_25.INIT0 = 16'h5999;
    defparam sub_1721_add_2_25.INIT1 = 16'h5999;
    defparam sub_1721_add_2_25.INJECT1_0 = "NO";
    defparam sub_1721_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27436), .COUT(n27437));
    defparam sub_1721_add_2_23.INIT0 = 16'h5999;
    defparam sub_1721_add_2_23.INIT1 = 16'h5999;
    defparam sub_1721_add_2_23.INJECT1_0 = "NO";
    defparam sub_1721_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27435), .COUT(n27436));
    defparam sub_1721_add_2_21.INIT0 = 16'h5999;
    defparam sub_1721_add_2_21.INIT1 = 16'h5999;
    defparam sub_1721_add_2_21.INJECT1_0 = "NO";
    defparam sub_1721_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27434), .COUT(n27435));
    defparam sub_1721_add_2_19.INIT0 = 16'h5999;
    defparam sub_1721_add_2_19.INIT1 = 16'h5999;
    defparam sub_1721_add_2_19.INJECT1_0 = "NO";
    defparam sub_1721_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27433), .COUT(n27434));
    defparam sub_1721_add_2_17.INIT0 = 16'h5999;
    defparam sub_1721_add_2_17.INIT1 = 16'h5999;
    defparam sub_1721_add_2_17.INJECT1_0 = "NO";
    defparam sub_1721_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27432), .COUT(n27433));
    defparam sub_1721_add_2_15.INIT0 = 16'h5999;
    defparam sub_1721_add_2_15.INIT1 = 16'h5999;
    defparam sub_1721_add_2_15.INJECT1_0 = "NO";
    defparam sub_1721_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27431), .COUT(n27432));
    defparam sub_1721_add_2_13.INIT0 = 16'h5999;
    defparam sub_1721_add_2_13.INIT1 = 16'h5999;
    defparam sub_1721_add_2_13.INJECT1_0 = "NO";
    defparam sub_1721_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27430), .COUT(n27431));
    defparam sub_1721_add_2_11.INIT0 = 16'h5999;
    defparam sub_1721_add_2_11.INIT1 = 16'h5999;
    defparam sub_1721_add_2_11.INJECT1_0 = "NO";
    defparam sub_1721_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27429), .COUT(n27430));
    defparam sub_1721_add_2_9.INIT0 = 16'h5999;
    defparam sub_1721_add_2_9.INIT1 = 16'h5999;
    defparam sub_1721_add_2_9.INJECT1_0 = "NO";
    defparam sub_1721_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27428), .COUT(n27429));
    defparam sub_1721_add_2_7.INIT0 = 16'h5999;
    defparam sub_1721_add_2_7.INIT1 = 16'h5999;
    defparam sub_1721_add_2_7.INJECT1_0 = "NO";
    defparam sub_1721_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27427), .COUT(n27428));
    defparam sub_1721_add_2_5.INIT0 = 16'h5999;
    defparam sub_1721_add_2_5.INIT1 = 16'h5999;
    defparam sub_1721_add_2_5.INJECT1_0 = "NO";
    defparam sub_1721_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27426), .COUT(n27427));
    defparam sub_1721_add_2_3.INIT0 = 16'h5999;
    defparam sub_1721_add_2_3.INIT1 = 16'h5999;
    defparam sub_1721_add_2_3.INJECT1_0 = "NO";
    defparam sub_1721_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1721_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27426));
    defparam sub_1721_add_2_1.INIT0 = 16'h0000;
    defparam sub_1721_add_2_1.INIT1 = 16'h5999;
    defparam sub_1721_add_2_1.INJECT1_0 = "NO";
    defparam sub_1721_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27425), .S1(n6986));
    defparam sub_1722_add_2_33.INIT0 = 16'hf555;
    defparam sub_1722_add_2_33.INIT1 = 16'h0000;
    defparam sub_1722_add_2_33.INJECT1_0 = "NO";
    defparam sub_1722_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27424), .COUT(n27425));
    defparam sub_1722_add_2_31.INIT0 = 16'hf555;
    defparam sub_1722_add_2_31.INIT1 = 16'hf555;
    defparam sub_1722_add_2_31.INJECT1_0 = "NO";
    defparam sub_1722_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27423), .COUT(n27424));
    defparam sub_1722_add_2_29.INIT0 = 16'hf555;
    defparam sub_1722_add_2_29.INIT1 = 16'hf555;
    defparam sub_1722_add_2_29.INJECT1_0 = "NO";
    defparam sub_1722_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27422), .COUT(n27423));
    defparam sub_1722_add_2_27.INIT0 = 16'hf555;
    defparam sub_1722_add_2_27.INIT1 = 16'hf555;
    defparam sub_1722_add_2_27.INJECT1_0 = "NO";
    defparam sub_1722_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27421), .COUT(n27422));
    defparam sub_1722_add_2_25.INIT0 = 16'hf555;
    defparam sub_1722_add_2_25.INIT1 = 16'hf555;
    defparam sub_1722_add_2_25.INJECT1_0 = "NO";
    defparam sub_1722_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27420), .COUT(n27421));
    defparam sub_1722_add_2_23.INIT0 = 16'hf555;
    defparam sub_1722_add_2_23.INIT1 = 16'hf555;
    defparam sub_1722_add_2_23.INJECT1_0 = "NO";
    defparam sub_1722_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27419), .COUT(n27420));
    defparam sub_1722_add_2_21.INIT0 = 16'hf555;
    defparam sub_1722_add_2_21.INIT1 = 16'hf555;
    defparam sub_1722_add_2_21.INJECT1_0 = "NO";
    defparam sub_1722_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27418), .COUT(n27419));
    defparam sub_1722_add_2_19.INIT0 = 16'hf555;
    defparam sub_1722_add_2_19.INIT1 = 16'hf555;
    defparam sub_1722_add_2_19.INJECT1_0 = "NO";
    defparam sub_1722_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27417), .COUT(n27418));
    defparam sub_1722_add_2_17.INIT0 = 16'hf555;
    defparam sub_1722_add_2_17.INIT1 = 16'hf555;
    defparam sub_1722_add_2_17.INJECT1_0 = "NO";
    defparam sub_1722_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27416), .COUT(n27417));
    defparam sub_1722_add_2_15.INIT0 = 16'hf555;
    defparam sub_1722_add_2_15.INIT1 = 16'hf555;
    defparam sub_1722_add_2_15.INJECT1_0 = "NO";
    defparam sub_1722_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27415), .COUT(n27416));
    defparam sub_1722_add_2_13.INIT0 = 16'hf555;
    defparam sub_1722_add_2_13.INIT1 = 16'hf555;
    defparam sub_1722_add_2_13.INJECT1_0 = "NO";
    defparam sub_1722_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27414), .COUT(n27415));
    defparam sub_1722_add_2_11.INIT0 = 16'hf555;
    defparam sub_1722_add_2_11.INIT1 = 16'hf555;
    defparam sub_1722_add_2_11.INJECT1_0 = "NO";
    defparam sub_1722_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27413), .COUT(n27414));
    defparam sub_1722_add_2_9.INIT0 = 16'hf555;
    defparam sub_1722_add_2_9.INIT1 = 16'hf555;
    defparam sub_1722_add_2_9.INJECT1_0 = "NO";
    defparam sub_1722_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27412), .COUT(n27413));
    defparam sub_1722_add_2_7.INIT0 = 16'hf555;
    defparam sub_1722_add_2_7.INIT1 = 16'hf555;
    defparam sub_1722_add_2_7.INJECT1_0 = "NO";
    defparam sub_1722_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27411), .COUT(n27412));
    defparam sub_1722_add_2_5.INIT0 = 16'hf555;
    defparam sub_1722_add_2_5.INIT1 = 16'hf555;
    defparam sub_1722_add_2_5.INJECT1_0 = "NO";
    defparam sub_1722_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27410), .COUT(n27411));
    defparam sub_1722_add_2_3.INIT0 = 16'hf555;
    defparam sub_1722_add_2_3.INIT1 = 16'hf555;
    defparam sub_1722_add_2_3.INJECT1_0 = "NO";
    defparam sub_1722_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1722_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27410));
    defparam sub_1722_add_2_1.INIT0 = 16'h0000;
    defparam sub_1722_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1722_add_2_1.INJECT1_0 = "NO";
    defparam sub_1722_add_2_1.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27877), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_33.INIT1 = 16'h0000;
    defparam count_2177_add_4_33.INJECT1_0 = "NO";
    defparam count_2177_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27876), .COUT(n27877), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_31.INJECT1_0 = "NO";
    defparam count_2177_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27875), .COUT(n27876), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_29.INJECT1_0 = "NO";
    defparam count_2177_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27874), .COUT(n27875), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_27.INJECT1_0 = "NO";
    defparam count_2177_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27873), .COUT(n27874), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_25.INJECT1_0 = "NO";
    defparam count_2177_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27872), .COUT(n27873), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_23.INJECT1_0 = "NO";
    defparam count_2177_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27871), .COUT(n27872), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_21.INJECT1_0 = "NO";
    defparam count_2177_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27870), .COUT(n27871), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_19.INJECT1_0 = "NO";
    defparam count_2177_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27869), .COUT(n27870), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_17.INJECT1_0 = "NO";
    defparam count_2177_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27868), .COUT(n27869), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_15.INJECT1_0 = "NO";
    defparam count_2177_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27867), .COUT(n27868), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_13.INJECT1_0 = "NO";
    defparam count_2177_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27866), .COUT(n27867), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_11.INJECT1_0 = "NO";
    defparam count_2177_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27865), .COUT(n27866), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_9.INJECT1_0 = "NO";
    defparam count_2177_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27864), .COUT(n27865), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_7.INJECT1_0 = "NO";
    defparam count_2177_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27863), .COUT(n27864), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_5.INJECT1_0 = "NO";
    defparam count_2177_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27862), .COUT(n27863), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2177_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2177_add_4_3.INJECT1_0 = "NO";
    defparam count_2177_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2177_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27862), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2177_add_4_1.INIT0 = 16'hF000;
    defparam count_2177_add_4_1.INIT1 = 16'h0555;
    defparam count_2177_add_4_1.INJECT1_0 = "NO";
    defparam count_2177_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module RCPeripheral
//

module RCPeripheral (\read_value[13] , n1, n32472, \read_value[13]_adj_43 , 
            read_value, n32375, n52, \register_addr[0] , databus_out, 
            n2, rw, databus, \read_value[12]_adj_45 , n1_adj_46, n4, 
            \read_value[12]_adj_47 , n2_adj_48, \read_value[11]_adj_49 , 
            n1_adj_50, \read_value[11]_adj_51 , \select[7] , n32504, 
            n32481, \register_addr[1] , n30427, n30283, n30284, n32505, 
            n30631, n29663, n11883, n30710, n30411, n2_adj_52, \read_value[10]_adj_53 , 
            n1_adj_54, \read_value[10]_adj_55 , \register_addr[4] , \read_size[0] , 
            \read_size[0]_adj_56 , \register_addr[5] , \read_size[0]_adj_57 , 
            \read_size[0]_adj_58 , n2_adj_59, n2_adj_60, \read_value[18]_adj_61 , 
            n1_adj_62, \read_value[18]_adj_63 , \read_value[2]_adj_64 , 
            n32374, \read_value[24]_adj_65 , n1_adj_66, n2_adj_67, \read_value[2]_adj_68 , 
            \read_value[2]_adj_69 , n32376, \read_value[9]_adj_70 , n1_adj_71, 
            \read_value[24]_adj_72 , \read_value[9]_adj_73 , n32455, \register_addr[2] , 
            \register_addr[3] , n30401, read_value_adj_186, n64, n2_adj_82, 
            \read_value[17]_adj_83 , n1_adj_84, \read_value[17]_adj_85 , 
            n2_adj_86, n2_adj_87, \read_value[16]_adj_88 , n1_adj_89, 
            \read_value[16]_adj_90 , read_size, \select[1] , n32486, 
            \sendcount[1] , n11271, n2_adj_92, \read_value[15]_adj_93 , 
            n1_adj_94, n2_adj_95, \read_value[15]_adj_96 , \read_value[23]_adj_97 , 
            n1_adj_98, n32381, n30423, n32345, \read_value[8]_adj_99 , 
            n1_adj_100, n1_adj_101, n2_adj_102, \read_value[14]_adj_103 , 
            n1_adj_104, \read_value[8]_adj_105 , \read_value[14]_adj_106 , 
            \read_value[1]_adj_107 , n6, \read_value[23]_adj_108 , n2_adj_109, 
            \read_value[1]_adj_110 , n2_adj_111, \read_value[22]_adj_112 , 
            n1_adj_113, \read_value[22]_adj_114 , n2_adj_115, n2_adj_116, 
            \read_value[30]_adj_117 , n1_adj_118, \read_value[19]_adj_119 , 
            n1_adj_120, n4_adj_121, \read_value[7]_adj_122 , \read_value[30]_adj_123 , 
            n2_adj_124, \read_value[19]_adj_125 , \read_size[2]_adj_126 , 
            \read_size[2]_adj_127 , \read_size[2]_adj_128 , \read_size[2]_adj_129 , 
            \read_value[7]_adj_130 , \read_value[7]_adj_131 , n34317, 
            \read_value[29]_adj_132 , n1_adj_133, n2_adj_134, n4_adj_135, 
            \read_value[6]_adj_136 , \read_value[6]_adj_137 , \read_value[6]_adj_138 , 
            \read_value[29]_adj_139 , n4_adj_140, \read_value[0]_adj_141 , 
            \read_value[0]_adj_142 , \read_value[0]_adj_143 , \read_value[21]_adj_144 , 
            n1_adj_145, n4_adj_146, \read_value[5]_adj_147 , \read_value[5]_adj_148 , 
            \read_value[5]_adj_149 , \read_value[21]_adj_150 , n2_adj_151, 
            \select[2] , \read_size[0]_adj_152 , n5, n32439, n6_adj_153, 
            n2_adj_154, \read_value[31]_adj_155 , n1_adj_156, \read_value[31]_adj_157 , 
            \reg_size[2] , n2_adj_158, \read_value[28]_adj_159 , n1_adj_160, 
            \read_value[28]_adj_161 , \read_value[20]_adj_162 , n1_adj_163, 
            n4_adj_164, \read_value[4]_adj_165 , \read_value[4]_adj_166 , 
            \read_value[4]_adj_167 , \read_value[20]_adj_168 , n2_adj_169, 
            \read_value[27]_adj_170 , n1_adj_171, \read_value[27]_adj_172 , 
            n2_adj_173, \read_value[26]_adj_174 , n1_adj_175, \read_value[26]_adj_176 , 
            n4_adj_177, \read_value[3]_adj_178 , \read_value[3]_adj_179 , 
            \read_value[3]_adj_180 , n2_adj_181, \read_value[25]_adj_182 , 
            n1_adj_183, \read_value[25]_adj_184 , debug_c_c, n28324, 
            GND_net, n32341, rc_ch8_c, n31024, n30913, n12030, n31005, 
            n28308, rc_ch7_c, n30995, n12031, n30929, rc_ch4_c, 
            n28304, n12138, n31000, n30969, n28317, rc_ch3_c, n1000, 
            n988, n32336, n14446, rc_ch2_c, n54, n4_adj_185, n12841, 
            n31049, n28312, rc_ch1_c, n30911) /* synthesis syn_module_defined=1 */ ;
    input \read_value[13] ;
    input n1;
    input n32472;
    input \read_value[13]_adj_43 ;
    input [31:0]read_value;
    input n32375;
    input n52;
    input \register_addr[0] ;
    input [31:0]databus_out;
    input n2;
    input rw;
    output [31:0]databus;
    input \read_value[12]_adj_45 ;
    input n1_adj_46;
    input n4;
    input \read_value[12]_adj_47 ;
    input n2_adj_48;
    input \read_value[11]_adj_49 ;
    input n1_adj_50;
    input \read_value[11]_adj_51 ;
    input \select[7] ;
    input n32504;
    input n32481;
    input \register_addr[1] ;
    output n30427;
    output n30283;
    output n30284;
    input n32505;
    output n30631;
    output n29663;
    input n11883;
    output n30710;
    output n30411;
    input n2_adj_52;
    input \read_value[10]_adj_53 ;
    input n1_adj_54;
    input \read_value[10]_adj_55 ;
    input \register_addr[4] ;
    input \read_size[0] ;
    input \read_size[0]_adj_56 ;
    input \register_addr[5] ;
    input \read_size[0]_adj_57 ;
    input \read_size[0]_adj_58 ;
    input n2_adj_59;
    input n2_adj_60;
    input \read_value[18]_adj_61 ;
    input n1_adj_62;
    input \read_value[18]_adj_63 ;
    input \read_value[2]_adj_64 ;
    input n32374;
    input \read_value[24]_adj_65 ;
    input n1_adj_66;
    input n2_adj_67;
    input \read_value[2]_adj_68 ;
    input \read_value[2]_adj_69 ;
    input n32376;
    input \read_value[9]_adj_70 ;
    input n1_adj_71;
    input \read_value[24]_adj_72 ;
    input \read_value[9]_adj_73 ;
    input n32455;
    input \register_addr[2] ;
    input \register_addr[3] ;
    output n30401;
    input [7:0]read_value_adj_186;
    input n64;
    input n2_adj_82;
    input \read_value[17]_adj_83 ;
    input n1_adj_84;
    input \read_value[17]_adj_85 ;
    input n2_adj_86;
    input n2_adj_87;
    input \read_value[16]_adj_88 ;
    input n1_adj_89;
    input \read_value[16]_adj_90 ;
    input [2:0]read_size;
    input \select[1] ;
    output n32486;
    input \sendcount[1] ;
    output n11271;
    input n2_adj_92;
    input \read_value[15]_adj_93 ;
    input n1_adj_94;
    input n2_adj_95;
    input \read_value[15]_adj_96 ;
    input \read_value[23]_adj_97 ;
    input n1_adj_98;
    input n32381;
    input n30423;
    output n32345;
    input \read_value[8]_adj_99 ;
    input n1_adj_100;
    input n1_adj_101;
    input n2_adj_102;
    input \read_value[14]_adj_103 ;
    input n1_adj_104;
    input \read_value[8]_adj_105 ;
    input \read_value[14]_adj_106 ;
    input \read_value[1]_adj_107 ;
    input n6;
    input \read_value[23]_adj_108 ;
    input n2_adj_109;
    input \read_value[1]_adj_110 ;
    input n2_adj_111;
    input \read_value[22]_adj_112 ;
    input n1_adj_113;
    input \read_value[22]_adj_114 ;
    input n2_adj_115;
    input n2_adj_116;
    input \read_value[30]_adj_117 ;
    input n1_adj_118;
    input \read_value[19]_adj_119 ;
    input n1_adj_120;
    input n4_adj_121;
    input \read_value[7]_adj_122 ;
    input \read_value[30]_adj_123 ;
    input n2_adj_124;
    input \read_value[19]_adj_125 ;
    input \read_size[2]_adj_126 ;
    input \read_size[2]_adj_127 ;
    input \read_size[2]_adj_128 ;
    input \read_size[2]_adj_129 ;
    input \read_value[7]_adj_130 ;
    input \read_value[7]_adj_131 ;
    input n34317;
    input \read_value[29]_adj_132 ;
    input n1_adj_133;
    input n2_adj_134;
    input n4_adj_135;
    input \read_value[6]_adj_136 ;
    input \read_value[6]_adj_137 ;
    input \read_value[6]_adj_138 ;
    input \read_value[29]_adj_139 ;
    input n4_adj_140;
    input \read_value[0]_adj_141 ;
    input \read_value[0]_adj_142 ;
    input \read_value[0]_adj_143 ;
    input \read_value[21]_adj_144 ;
    input n1_adj_145;
    input n4_adj_146;
    input \read_value[5]_adj_147 ;
    input \read_value[5]_adj_148 ;
    input \read_value[5]_adj_149 ;
    input \read_value[21]_adj_150 ;
    input n2_adj_151;
    input \select[2] ;
    input \read_size[0]_adj_152 ;
    output n5;
    input n32439;
    output n6_adj_153;
    input n2_adj_154;
    input \read_value[31]_adj_155 ;
    input n1_adj_156;
    input \read_value[31]_adj_157 ;
    output \reg_size[2] ;
    input n2_adj_158;
    input \read_value[28]_adj_159 ;
    input n1_adj_160;
    input \read_value[28]_adj_161 ;
    input \read_value[20]_adj_162 ;
    input n1_adj_163;
    input n4_adj_164;
    input \read_value[4]_adj_165 ;
    input \read_value[4]_adj_166 ;
    input \read_value[4]_adj_167 ;
    input \read_value[20]_adj_168 ;
    input n2_adj_169;
    input \read_value[27]_adj_170 ;
    input n1_adj_171;
    input \read_value[27]_adj_172 ;
    input n2_adj_173;
    input \read_value[26]_adj_174 ;
    input n1_adj_175;
    input \read_value[26]_adj_176 ;
    input n4_adj_177;
    input \read_value[3]_adj_178 ;
    input \read_value[3]_adj_179 ;
    input \read_value[3]_adj_180 ;
    input n2_adj_181;
    input \read_value[25]_adj_182 ;
    input n1_adj_183;
    input \read_value[25]_adj_184 ;
    input debug_c_c;
    input n28324;
    input GND_net;
    input n32341;
    input rc_ch8_c;
    output n31024;
    output n30913;
    input n12030;
    output n31005;
    input n28308;
    input rc_ch7_c;
    output n30995;
    input n12031;
    output n30929;
    input rc_ch4_c;
    input n28304;
    input n12138;
    output n31000;
    output n30969;
    input n28317;
    input rc_ch3_c;
    output n1000;
    output n988;
    input n32336;
    input n14446;
    input rc_ch2_c;
    output n54;
    output n4_adj_185;
    input n12841;
    output n31049;
    input n28312;
    input rc_ch1_c;
    output n30911;
    
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n8, n10;
    wire [7:0]\register[6] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    
    wire n31516, n10_adj_137, n8_adj_138, n32185;
    wire [7:0]\register[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    wire [7:0]\register[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    
    wire n31519, n1054;
    wire [7:0]\register[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    
    wire n31520, n13, n12, n6_c;
    wire [7:0]\register[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    wire [7:0]\register[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(209[13:21])
    
    wire n32186, n32188, n994, n32189, n32222, n10_adj_142, n8_adj_144, 
        n32219;
    wire [2:0]read_size_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(213[12:21])
    
    wire n176, n979, n32223, n32220, n10_adj_148, n8_adj_150, n19, 
        n22, n25, n31900, n32258, n18, n21, n24, n32259, n32473;
    wire [7:0]read_value_adj_368;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(212[12:22])
    
    wire n7, n7_adj_158, n7_adj_159, n7_adj_160, n31485, n7_adj_161, 
        n7_adj_162, n7_adj_163, n10_adj_164, n10_adj_166, n8_adj_168, 
        n10_adj_173, n8_adj_174, n10_adj_176, n32256, n32255, n8_adj_180, 
        n32431, n32273, n32274, n32276, n10_adj_188, n8_adj_190, 
        n31897, n1039, n32277, n10_adj_194, n10_adj_196, n8_adj_198, 
        n31898, n31901, n10_adj_202, n8_adj_204, n10_adj_206, n8_adj_210, 
        n8_adj_212, n14, n10_adj_215, n7_adj_216, n1009, n32106, 
        n10_adj_217, n8_adj_219, n12_adj_225, n32225, n32105, n32103, 
        n32102, n31517, n31522, n32279, n31903, n32261, n31491, 
        n32108, n10_adj_234, n32191, n8_adj_236, n10_adj_240, n10_adj_242, 
        n8_adj_244, n8_adj_246, n32278, n32275, n13_adj_248, n12_adj_250, 
        n6_adj_251, n10_adj_253, n31488, n1024, n31489, n32260, 
        n32257, n10_adj_256, n8_adj_265, n10_adj_269, n13_adj_271, 
        n12_adj_273, n6_adj_274, n10_adj_276, n13_adj_283, n12_adj_285, 
        n6_adj_286, n32224, n32221, n31486, n10_adj_288, n8_adj_291, 
        n13_adj_295, n12_adj_297, n6_adj_298, n10_adj_300, n32190, 
        n32187, n31487, n31521, n31518, n10_adj_307, n10_adj_312, 
        n8_adj_314, n10_adj_319, n8_adj_321, n32107, n32104, n8_adj_325, 
        n13_adj_327, n12_adj_329, n6_adj_330, n10_adj_332, n10_adj_339, 
        n31902, n31899, n31490, n8_adj_341, n10_adj_345, n8_adj_347, 
        n13_adj_351, n12_adj_353, n6_adj_354, n10_adj_356, n10_adj_359, 
        n8_adj_363;
    
    LUT4 i4_4_lut (.A(\read_value[13] ), .B(n8), .C(n1), .D(n32472), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut.init = 16'hfefc;
    LUT4 i2_4_lut (.A(\read_value[13]_adj_43 ), .B(read_value[13]), .C(n32375), 
         .D(n52), .Z(n8)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_24979 (.A(\register[6] [7]), .B(\register_addr[0] ), 
         .Z(n31516)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_24979.init = 16'h2222;
    LUT4 i5_4_lut (.A(databus_out[12]), .B(n10_adj_137), .C(n2), .D(rw), 
         .Z(databus[12])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_264 (.A(\read_value[12]_adj_45 ), .B(n8_adj_138), 
         .C(n1_adj_46), .D(n32472), .Z(n10_adj_137)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_264.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_25180 (.A(\register[6] [1]), .B(\register_addr[0] ), 
         .Z(n32185)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_25180.init = 16'h2222;
    LUT4 n1054_bdd_3_lut_24935 (.A(\register[2] [7]), .B(\register[3] [7]), 
         .C(\register_addr[0] ), .Z(n31519)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1054_bdd_3_lut_24935.init = 16'hcaca;
    LUT4 n1054_bdd_3_lut_25157 (.A(n1054), .B(\register_addr[0] ), .C(\register[1] [7]), 
         .Z(n31520)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1054_bdd_3_lut_25157.init = 16'he2e2;
    LUT4 i7_4_lut (.A(n13), .B(n4), .C(n12), .D(n6_c), .Z(databus[2])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 register_addr_1__bdd_3_lut_25181 (.A(\register_addr[0] ), .B(\register[4] [1]), 
         .C(\register[5] [1]), .Z(n32186)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_25181.init = 16'he4e4;
    LUT4 n994_bdd_3_lut_25175 (.A(\register[2] [1]), .B(\register[3] [1]), 
         .C(\register_addr[0] ), .Z(n32188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n994_bdd_3_lut_25175.init = 16'hcaca;
    LUT4 i2_4_lut_adj_265 (.A(\read_value[12]_adj_47 ), .B(read_value[12]), 
         .C(n32375), .D(n52), .Z(n8_adj_138)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_265.init = 16'heca0;
    LUT4 n994_bdd_3_lut_25977 (.A(n994), .B(\register_addr[0] ), .C(\register[1] [1]), 
         .Z(n32189)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n994_bdd_3_lut_25977.init = 16'he2e2;
    LUT4 n979_bdd_3_lut_25186 (.A(\register[2] [0]), .B(\register[3] [0]), 
         .C(\register_addr[0] ), .Z(n32222)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n979_bdd_3_lut_25186.init = 16'hcaca;
    LUT4 i5_4_lut_adj_266 (.A(databus_out[11]), .B(n10_adj_142), .C(n2_adj_48), 
         .D(rw), .Z(databus[11])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_266.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_267 (.A(\read_value[11]_adj_49 ), .B(n8_adj_144), 
         .C(n1_adj_50), .D(n32472), .Z(n10_adj_142)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_267.init = 16'hfefc;
    LUT4 i2_4_lut_adj_268 (.A(\read_value[11]_adj_51 ), .B(read_value[11]), 
         .C(n32375), .D(n52), .Z(n8_adj_144)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_268.init = 16'heca0;
    LUT4 register_addr_1__bdd_2_lut_25203 (.A(\register[6] [0]), .B(\register_addr[0] ), 
         .Z(n32219)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_25203.init = 16'h2222;
    FD1S3AX read_size_i1 (.D(n176), .CK(\select[7] ), .Q(read_size_c[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_size_i1.GSR = "ENABLED";
    LUT4 n979_bdd_3_lut_25900 (.A(n979), .B(\register_addr[0] ), .C(\register[1] [0]), 
         .Z(n32223)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n979_bdd_3_lut_25900.init = 16'he2e2;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32504), .B(n32481), .C(\register_addr[1] ), 
         .D(n30427), .Z(n30283)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_4_lut_adj_269 (.A(n32504), .B(n32481), .C(\register_addr[1] ), 
         .D(n30427), .Z(n30284)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_269.init = 16'h1000;
    LUT4 i24802_2_lut_3_lut_4_lut (.A(n32504), .B(n32481), .C(\register_addr[1] ), 
         .D(n32505), .Z(n30631)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i24802_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_4_lut_adj_270 (.A(n32504), .B(n32481), .C(\register_addr[1] ), 
         .D(n32505), .Z(n29663)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_270.init = 16'h0010;
    LUT4 register_addr_1__bdd_3_lut_25204 (.A(\register_addr[0] ), .B(\register[4] [0]), 
         .C(\register[5] [0]), .Z(n32220)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_25204.init = 16'he4e4;
    LUT4 i24741_2_lut_3_lut_4_lut (.A(n32504), .B(n32481), .C(\register_addr[1] ), 
         .D(n11883), .Z(n30710)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i24741_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_4_lut_adj_271 (.A(n32504), .B(n32481), .C(\register_addr[1] ), 
         .D(n11883), .Z(n30411)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_271.init = 16'h0010;
    LUT4 i5_4_lut_adj_272 (.A(databus_out[10]), .B(n10_adj_148), .C(n2_adj_52), 
         .D(rw), .Z(databus[10])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_272.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_273 (.A(\read_value[10]_adj_53 ), .B(n8_adj_150), 
         .C(n1_adj_54), .D(n32472), .Z(n10_adj_148)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_273.init = 16'hfefc;
    LUT4 i2_4_lut_adj_274 (.A(\read_value[10]_adj_55 ), .B(read_value[10]), 
         .C(n32375), .D(n52), .Z(n8_adj_150)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_274.init = 16'heca0;
    PFUMX i38 (.BLUT(n19), .ALUT(n22), .C0(\register_addr[4] ), .Z(n25));
    LUT4 i24540_3_lut (.A(\read_size[0] ), .B(\read_size[0]_adj_56 ), .C(\register_addr[5] ), 
         .Z(n19)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24540_3_lut.init = 16'hcaca;
    LUT4 i24541_3_lut (.A(\read_size[0]_adj_57 ), .B(\read_size[0]_adj_58 ), 
         .C(\register_addr[5] ), .Z(n22)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24541_3_lut.init = 16'hcaca;
    LUT4 \register_1[[5__bdd_3_lut_25193  (.A(\register[2] [5]), .B(\register[3] [5]), 
         .C(\register_addr[0] ), .Z(n31900)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[5__bdd_3_lut_25193 .init = 16'hcaca;
    LUT4 \register_1[[4__bdd_3_lut_25853  (.A(\register[2] [4]), .B(\register[3] [4]), 
         .C(\register_addr[0] ), .Z(n32258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \register_1[[4__bdd_3_lut_25853 .init = 16'hcaca;
    PFUMX i37 (.BLUT(n18), .ALUT(n21), .C0(\register_addr[4] ), .Z(n24));
    LUT4 \register_1[[4__bdd_2_lut_25854  (.A(\register[1] [4]), .B(\register_addr[0] ), 
         .Z(n32259)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[4__bdd_2_lut_25854 .init = 16'h8888;
    LUT4 i14_2_lut_rep_379 (.A(\select[7] ), .B(rw), .Z(n32473)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam i14_2_lut_rep_379.init = 16'h8888;
    LUT4 Select_3619_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_368[6]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3619_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3620_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_368[5]), 
         .Z(n7_adj_158)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3620_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3618_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_368[7]), 
         .Z(n7_adj_159)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3618_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3625_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_368[0]), 
         .Z(n7_adj_160)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3625_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 register_addr_1__bdd_2_lut_24926 (.A(\register[6] [3]), .B(\register_addr[0] ), 
         .Z(n31485)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_24926.init = 16'h2222;
    LUT4 Select_3623_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_368[2]), 
         .Z(n7_adj_161)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3623_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3622_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_368[3]), 
         .Z(n7_adj_162)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3622_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 Select_3621_i7_2_lut_3_lut (.A(\select[7] ), .B(rw), .C(read_value_adj_368[4]), 
         .Z(n7_adj_163)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(216[19:32])
    defparam Select_3621_i7_2_lut_3_lut.init = 16'h8080;
    LUT4 i5_4_lut_adj_275 (.A(databus_out[18]), .B(n10_adj_164), .C(n2_adj_59), 
         .D(rw), .Z(databus[18])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_275.init = 16'hfcfe;
    LUT4 i5_4_lut_adj_276 (.A(databus_out[24]), .B(n10_adj_166), .C(n2_adj_60), 
         .D(rw), .Z(databus[24])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_276.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_277 (.A(\read_value[18]_adj_61 ), .B(n8_adj_168), 
         .C(n1_adj_62), .D(n32472), .Z(n10_adj_164)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_277.init = 16'hfefc;
    LUT4 i2_4_lut_adj_278 (.A(\read_value[18]_adj_63 ), .B(read_value[18]), 
         .C(n32375), .D(n52), .Z(n8_adj_168)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_278.init = 16'heca0;
    LUT4 i5_4_lut_adj_279 (.A(\read_value[2]_adj_64 ), .B(n10_adj_173), 
         .C(n7_adj_161), .D(n32374), .Z(n13)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_279.init = 16'hfefc;
    LUT4 i4_4_lut_adj_280 (.A(\read_value[24]_adj_65 ), .B(n8_adj_174), 
         .C(n1_adj_66), .D(n32472), .Z(n10_adj_166)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_280.init = 16'hfefc;
    LUT4 i5_4_lut_adj_281 (.A(databus_out[9]), .B(n10_adj_176), .C(n2_adj_67), 
         .D(rw), .Z(databus[9])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_281.init = 16'hfcfe;
    LUT4 register_addr_1__bdd_3_lut_25227 (.A(\register_addr[0] ), .B(\register[4] [4]), 
         .C(\register[5] [4]), .Z(n32256)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_25227.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_25226 (.A(\register[6] [4]), .B(\register_addr[0] ), 
         .Z(n32255)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_25226.init = 16'h2222;
    LUT4 i4_4_lut_adj_282 (.A(\read_value[2]_adj_68 ), .B(\read_value[2]_adj_69 ), 
         .C(n32376), .D(n32472), .Z(n12)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_282.init = 16'heca0;
    LUT4 i4_4_lut_adj_283 (.A(\read_value[9]_adj_70 ), .B(n8_adj_180), .C(n1_adj_71), 
         .D(n32472), .Z(n10_adj_176)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_283.init = 16'hfefc;
    LUT4 i2_4_lut_adj_284 (.A(\read_value[24]_adj_72 ), .B(read_value[24]), 
         .C(n32375), .D(n52), .Z(n8_adj_174)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_284.init = 16'heca0;
    LUT4 i2_4_lut_adj_285 (.A(\read_value[9]_adj_73 ), .B(read_value[9]), 
         .C(n32375), .D(n52), .Z(n8_adj_180)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_285.init = 16'heca0;
    LUT4 i2_4_lut_rep_337 (.A(n32455), .B(\register_addr[2] ), .C(\register_addr[3] ), 
         .D(n30401), .Z(n32431)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(221[7:31])
    defparam i2_4_lut_rep_337.init = 16'hfefa;
    LUT4 i14560_1_lut_4_lut (.A(n32455), .B(\register_addr[2] ), .C(\register_addr[3] ), 
         .D(n30401), .Z(n176)) /* synthesis lut_function=(!(A+(B (C+(D))+!B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(221[7:31])
    defparam i14560_1_lut_4_lut.init = 16'h0105;
    LUT4 register_addr_1__bdd_2_lut (.A(\register[6] [6]), .B(\register_addr[0] ), 
         .Z(n32273)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut.init = 16'h2222;
    LUT4 register_addr_1__bdd_3_lut (.A(\register_addr[0] ), .B(\register[4] [6]), 
         .C(\register[5] [6]), .Z(n32274)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut.init = 16'he4e4;
    LUT4 n1039_bdd_3_lut_25230 (.A(\register[2] [6]), .B(\register[3] [6]), 
         .C(\register_addr[0] ), .Z(n32276)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1039_bdd_3_lut_25230.init = 16'hcaca;
    LUT4 Select_3623_i6_2_lut (.A(databus_out[2]), .B(rw), .Z(n6_c)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3623_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_286 (.A(read_value[2]), .B(read_value_adj_186[2]), 
         .C(n52), .D(n64), .Z(n10_adj_173)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_286.init = 16'heca0;
    LUT4 i5_4_lut_adj_287 (.A(databus_out[17]), .B(n10_adj_188), .C(n2_adj_82), 
         .D(rw), .Z(databus[17])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_287.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_288 (.A(\read_value[17]_adj_83 ), .B(n8_adj_190), 
         .C(n1_adj_84), .D(n32472), .Z(n10_adj_188)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_288.init = 16'hfefc;
    LUT4 register_addr_1__bdd_2_lut_25143 (.A(\register[6] [5]), .B(\register_addr[0] ), 
         .Z(n31897)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_25143.init = 16'h2222;
    LUT4 i2_4_lut_adj_289 (.A(\read_value[17]_adj_85 ), .B(read_value[17]), 
         .C(n32375), .D(n52), .Z(n8_adj_190)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_289.init = 16'heca0;
    LUT4 n1039_bdd_3_lut_25840 (.A(n1039), .B(\register_addr[0] ), .C(\register[1] [6]), 
         .Z(n32277)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1039_bdd_3_lut_25840.init = 16'he2e2;
    LUT4 i5_4_lut_adj_290 (.A(databus_out[23]), .B(n10_adj_194), .C(n2_adj_86), 
         .D(rw), .Z(databus[23])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_290.init = 16'hfcfe;
    LUT4 i5_4_lut_adj_291 (.A(databus_out[16]), .B(n10_adj_196), .C(n2_adj_87), 
         .D(rw), .Z(databus[16])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_291.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_292 (.A(\read_value[16]_adj_88 ), .B(n8_adj_198), 
         .C(n1_adj_89), .D(n32472), .Z(n10_adj_196)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_292.init = 16'hfefc;
    LUT4 i2_4_lut_adj_293 (.A(\read_value[16]_adj_90 ), .B(read_value[16]), 
         .C(n32375), .D(n52), .Z(n8_adj_198)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_293.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_25144 (.A(\register_addr[0] ), .B(\register[4] [5]), 
         .C(\register[5] [5]), .Z(n31898)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_25144.init = 16'he4e4;
    LUT4 Select_3633_i1_2_lut_rep_392 (.A(read_size[1]), .B(\select[1] ), 
         .Z(n32486)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_3633_i1_2_lut_rep_392.init = 16'h8888;
    LUT4 \register_1[[5__bdd_2_lut_25194  (.A(\register[1] [5]), .B(\register_addr[0] ), 
         .Z(n31901)) /* synthesis lut_function=(A (B)) */ ;
    defparam \register_1[[5__bdd_2_lut_25194 .init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(read_size[1]), .B(\select[1] ), .C(\sendcount[1] ), 
         .Z(n11271)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7878;
    LUT4 i5_4_lut_adj_294 (.A(databus_out[15]), .B(n10_adj_202), .C(n2_adj_92), 
         .D(rw), .Z(databus[15])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_294.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_295 (.A(\read_value[15]_adj_93 ), .B(n8_adj_204), 
         .C(n1_adj_94), .D(n32472), .Z(n10_adj_202)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_295.init = 16'hfefc;
    LUT4 i5_4_lut_adj_296 (.A(databus_out[8]), .B(n10_adj_206), .C(n2_adj_95), 
         .D(rw), .Z(databus[8])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_296.init = 16'hfcfe;
    LUT4 i2_4_lut_adj_297 (.A(\read_value[15]_adj_96 ), .B(read_value[15]), 
         .C(n32375), .D(n52), .Z(n8_adj_204)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_297.init = 16'heca0;
    LUT4 i4_4_lut_adj_298 (.A(\read_value[23]_adj_97 ), .B(n8_adj_210), 
         .C(n1_adj_98), .D(n32472), .Z(n10_adj_194)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_298.init = 16'hfefc;
    LUT4 i1_2_lut_rep_251_4_lut (.A(rw), .B(n30427), .C(n32381), .D(n30423), 
         .Z(n32345)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_rep_251_4_lut.init = 16'h4000;
    LUT4 i4_4_lut_adj_299 (.A(\read_value[8]_adj_99 ), .B(n8_adj_212), .C(n1_adj_100), 
         .D(n32472), .Z(n10_adj_206)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_299.init = 16'hfefc;
    LUT4 i7_4_lut_adj_300 (.A(n1_adj_101), .B(n14), .C(n10_adj_215), .D(n7_adj_216), 
         .Z(databus[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_300.init = 16'hfffe;
    LUT4 n1009_bdd_3_lut_25165 (.A(n1009), .B(\register_addr[0] ), .C(\register[1] [2]), 
         .Z(n32106)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1009_bdd_3_lut_25165.init = 16'he2e2;
    LUT4 i5_4_lut_adj_301 (.A(databus_out[14]), .B(n10_adj_217), .C(n2_adj_102), 
         .D(rw), .Z(databus[14])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_301.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_302 (.A(\read_value[14]_adj_103 ), .B(n8_adj_219), 
         .C(n1_adj_104), .D(n32472), .Z(n10_adj_217)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_302.init = 16'hfefc;
    LUT4 i2_4_lut_adj_303 (.A(\read_value[8]_adj_105 ), .B(read_value[8]), 
         .C(n32375), .D(n52), .Z(n8_adj_212)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_303.init = 16'heca0;
    LUT4 i2_4_lut_adj_304 (.A(\read_value[14]_adj_106 ), .B(read_value[14]), 
         .C(n32375), .D(n52), .Z(n8_adj_219)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_304.init = 16'heca0;
    LUT4 i6_4_lut (.A(\read_value[1]_adj_107 ), .B(n12_adj_225), .C(n6), 
         .D(n32375), .Z(n14)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut.init = 16'hfefc;
    FD1S3IX read_value__i0 (.D(n32225), .CK(\select[7] ), .CD(n32431), 
            .Q(read_value_adj_368[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 n1009_bdd_3_lut_25147 (.A(\register[2] [2]), .B(\register[3] [2]), 
         .C(\register_addr[0] ), .Z(n32105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1009_bdd_3_lut_25147.init = 16'hcaca;
    LUT4 register_addr_1__bdd_3_lut_25170 (.A(\register_addr[0] ), .B(\register[4] [2]), 
         .C(\register[5] [2]), .Z(n32103)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_25170.init = 16'he4e4;
    LUT4 register_addr_1__bdd_2_lut_25169 (.A(\register[6] [2]), .B(\register_addr[0] ), 
         .Z(n32102)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam register_addr_1__bdd_2_lut_25169.init = 16'h2222;
    LUT4 i2_4_lut_adj_305 (.A(read_value[1]), .B(read_value_adj_186[1]), 
         .C(n52), .D(n64), .Z(n10_adj_215)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_305.init = 16'heca0;
    LUT4 i2_4_lut_adj_306 (.A(\read_value[23]_adj_108 ), .B(read_value[23]), 
         .C(n32375), .D(n52), .Z(n8_adj_210)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_306.init = 16'heca0;
    LUT4 register_addr_1__bdd_3_lut_24980 (.A(\register_addr[0] ), .B(\register[4] [7]), 
         .C(\register[5] [7]), .Z(n31517)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_24980.init = 16'he4e4;
    LUT4 i5_4_lut_adj_307 (.A(databus_out[13]), .B(n10), .C(n2_adj_109), 
         .D(rw), .Z(databus[13])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_307.init = 16'hfcfe;
    LUT4 Select_3624_i7_2_lut (.A(databus_out[1]), .B(rw), .Z(n7_adj_216)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3624_i7_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_308 (.A(\read_value[1]_adj_110 ), .B(read_value_adj_368[1]), 
         .C(n32376), .D(n32473), .Z(n12_adj_225)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_308.init = 16'heca0;
    FD1S3IX read_value__i7 (.D(n31522), .CK(\select[7] ), .CD(n32431), 
            .Q(read_value_adj_368[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1S3IX read_value__i6 (.D(n32279), .CK(\select[7] ), .CD(n32431), 
            .Q(read_value_adj_368[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1S3IX read_value__i5 (.D(n31903), .CK(\select[7] ), .CD(n32431), 
            .Q(read_value_adj_368[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1S3IX read_value__i4 (.D(n32261), .CK(\select[7] ), .CD(n32431), 
            .Q(read_value_adj_368[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1S3IX read_value__i3 (.D(n31491), .CK(\select[7] ), .CD(n32431), 
            .Q(read_value_adj_368[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1S3IX read_value__i2 (.D(n32108), .CK(\select[7] ), .CD(n32431), 
            .Q(read_value_adj_368[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i2.GSR = "ENABLED";
    LUT4 i5_4_lut_adj_309 (.A(databus_out[22]), .B(n10_adj_234), .C(n2_adj_111), 
         .D(rw), .Z(databus[22])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_309.init = 16'hfcfe;
    FD1S3IX read_value__i1 (.D(n32191), .CK(\select[7] ), .CD(n32431), 
            .Q(read_value_adj_368[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=622, LSE_RLINE=634 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(219[9] 231[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i4_4_lut_adj_310 (.A(\read_value[22]_adj_112 ), .B(n8_adj_236), 
         .C(n1_adj_113), .D(n32472), .Z(n10_adj_234)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_310.init = 16'hfefc;
    LUT4 i2_4_lut_adj_311 (.A(\read_value[22]_adj_114 ), .B(read_value[22]), 
         .C(n32375), .D(n52), .Z(n8_adj_236)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_311.init = 16'heca0;
    LUT4 i5_4_lut_adj_312 (.A(databus_out[30]), .B(n10_adj_240), .C(n2_adj_115), 
         .D(rw), .Z(databus[30])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_312.init = 16'hfcfe;
    LUT4 i5_4_lut_adj_313 (.A(databus_out[19]), .B(n10_adj_242), .C(n2_adj_116), 
         .D(rw), .Z(databus[19])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_313.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_314 (.A(\read_value[30]_adj_117 ), .B(n8_adj_244), 
         .C(n1_adj_118), .D(n32472), .Z(n10_adj_240)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_314.init = 16'hfefc;
    LUT4 i4_4_lut_adj_315 (.A(\read_value[19]_adj_119 ), .B(n8_adj_246), 
         .C(n1_adj_120), .D(n32472), .Z(n10_adj_242)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_315.init = 16'hfefc;
    L6MUX21 i25233 (.D0(n32278), .D1(n32275), .SD(\register_addr[2] ), 
            .Z(n32279));
    PFUMX i25231 (.BLUT(n32277), .ALUT(n32276), .C0(\register_addr[1] ), 
          .Z(n32278));
    PFUMX i25228 (.BLUT(n32274), .ALUT(n32273), .C0(\register_addr[1] ), 
          .Z(n32275));
    LUT4 i7_4_lut_adj_316 (.A(n13_adj_248), .B(n4_adj_121), .C(n12_adj_250), 
         .D(n6_adj_251), .Z(databus[7])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_316.init = 16'hfffe;
    LUT4 i5_4_lut_adj_317 (.A(\read_value[7]_adj_122 ), .B(n10_adj_253), 
         .C(n7_adj_159), .D(n32374), .Z(n13_adj_248)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_317.init = 16'hfefc;
    LUT4 n1024_bdd_3_lut_24918 (.A(\register[2] [3]), .B(\register[3] [3]), 
         .C(\register_addr[0] ), .Z(n31488)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1024_bdd_3_lut_24918.init = 16'hcaca;
    LUT4 i2_4_lut_adj_318 (.A(\read_value[30]_adj_123 ), .B(read_value[30]), 
         .C(n32375), .D(n52), .Z(n8_adj_244)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_318.init = 16'heca0;
    LUT4 n1024_bdd_3_lut_25199 (.A(n1024), .B(\register_addr[0] ), .C(\register[1] [3]), 
         .Z(n31489)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n1024_bdd_3_lut_25199.init = 16'he2e2;
    L6MUX21 i25216 (.D0(n32260), .D1(n32257), .SD(\register_addr[2] ), 
            .Z(n32261));
    PFUMX i25214 (.BLUT(n32259), .ALUT(n32258), .C0(\register_addr[1] ), 
          .Z(n32260));
    PFUMX i25212 (.BLUT(n32256), .ALUT(n32255), .C0(\register_addr[1] ), 
          .Z(n32257));
    LUT4 i5_4_lut_adj_319 (.A(databus_out[29]), .B(n10_adj_256), .C(n2_adj_124), 
         .D(rw), .Z(databus[29])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_319.init = 16'hfcfe;
    LUT4 i2_4_lut_adj_320 (.A(\read_value[19]_adj_125 ), .B(read_value[19]), 
         .C(n32375), .D(n52), .Z(n8_adj_246)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_320.init = 16'heca0;
    LUT4 i39_3_lut (.A(\read_size[2]_adj_126 ), .B(\read_size[2]_adj_127 ), 
         .C(\register_addr[5] ), .Z(n18)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i39_3_lut.init = 16'hcaca;
    LUT4 i38_3_lut (.A(\read_size[2]_adj_128 ), .B(\read_size[2]_adj_129 ), 
         .C(\register_addr[5] ), .Z(n21)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38_3_lut.init = 16'hcaca;
    LUT4 i4_4_lut_adj_321 (.A(\read_value[7]_adj_130 ), .B(\read_value[7]_adj_131 ), 
         .C(n32376), .D(n32472), .Z(n12_adj_250)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_321.init = 16'heca0;
    LUT4 Select_3618_i6_2_lut (.A(databus_out[7]), .B(n34317), .Z(n6_adj_251)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3618_i6_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_322 (.A(\read_value[29]_adj_132 ), .B(n8_adj_265), 
         .C(n1_adj_133), .D(n32472), .Z(n10_adj_256)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_322.init = 16'hfefc;
    LUT4 i2_4_lut_adj_323 (.A(read_value[7]), .B(read_value_adj_186[7]), 
         .C(n52), .D(n64), .Z(n10_adj_253)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_323.init = 16'heca0;
    LUT4 i5_4_lut_adj_324 (.A(databus_out[21]), .B(n10_adj_269), .C(n2_adj_134), 
         .D(rw), .Z(databus[21])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_324.init = 16'hfcfe;
    LUT4 i7_4_lut_adj_325 (.A(n13_adj_271), .B(n4_adj_135), .C(n12_adj_273), 
         .D(n6_adj_274), .Z(databus[6])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_325.init = 16'hfffe;
    LUT4 i5_4_lut_adj_326 (.A(\read_value[6]_adj_136 ), .B(n10_adj_276), 
         .C(n7), .D(n32374), .Z(n13_adj_271)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_326.init = 16'hfefc;
    LUT4 i4_4_lut_adj_327 (.A(\read_value[6]_adj_137 ), .B(\read_value[6]_adj_138 ), 
         .C(n32376), .D(n32472), .Z(n12_adj_273)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_327.init = 16'heca0;
    LUT4 i2_4_lut_adj_328 (.A(\read_value[29]_adj_139 ), .B(read_value[29]), 
         .C(n32375), .D(n52), .Z(n8_adj_265)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_328.init = 16'heca0;
    LUT4 Select_3619_i6_2_lut (.A(databus_out[6]), .B(n34317), .Z(n6_adj_274)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3619_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_329 (.A(read_value[6]), .B(read_value_adj_186[6]), 
         .C(n52), .D(n64), .Z(n10_adj_276)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_329.init = 16'heca0;
    LUT4 i7_4_lut_adj_330 (.A(n13_adj_283), .B(n4_adj_140), .C(n12_adj_285), 
         .D(n6_adj_286), .Z(databus[0])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_330.init = 16'hfffe;
    L6MUX21 i25189 (.D0(n32224), .D1(n32221), .SD(\register_addr[2] ), 
            .Z(n32225));
    LUT4 register_addr_1__bdd_3_lut_24927 (.A(\register_addr[0] ), .B(\register[4] [3]), 
         .C(\register[5] [3]), .Z(n31486)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam register_addr_1__bdd_3_lut_24927.init = 16'he4e4;
    LUT4 i5_4_lut_adj_331 (.A(\read_value[0]_adj_141 ), .B(n10_adj_288), 
         .C(n7_adj_160), .D(n32374), .Z(n13_adj_283)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_331.init = 16'hfefc;
    LUT4 i4_4_lut_adj_332 (.A(\read_value[0]_adj_142 ), .B(\read_value[0]_adj_143 ), 
         .C(n32376), .D(n32472), .Z(n12_adj_285)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_332.init = 16'heca0;
    PFUMX i25187 (.BLUT(n32223), .ALUT(n32222), .C0(\register_addr[1] ), 
          .Z(n32224));
    LUT4 i4_4_lut_adj_333 (.A(\read_value[21]_adj_144 ), .B(n8_adj_291), 
         .C(n1_adj_145), .D(n32472), .Z(n10_adj_269)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_333.init = 16'hfefc;
    LUT4 Select_3625_i6_2_lut (.A(databus_out[0]), .B(n34317), .Z(n6_adj_286)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3625_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_334 (.A(read_value[0]), .B(read_value_adj_186[0]), 
         .C(n52), .D(n64), .Z(n10_adj_288)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_334.init = 16'heca0;
    LUT4 i7_4_lut_adj_335 (.A(n13_adj_295), .B(n4_adj_146), .C(n12_adj_297), 
         .D(n6_adj_298), .Z(databus[5])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_335.init = 16'hfffe;
    LUT4 i5_4_lut_adj_336 (.A(\read_value[5]_adj_147 ), .B(n10_adj_300), 
         .C(n7_adj_158), .D(n32374), .Z(n13_adj_295)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_336.init = 16'hfefc;
    LUT4 i4_4_lut_adj_337 (.A(\read_value[5]_adj_148 ), .B(\read_value[5]_adj_149 ), 
         .C(n32376), .D(n32472), .Z(n12_adj_297)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_337.init = 16'heca0;
    LUT4 Select_3620_i6_2_lut (.A(databus_out[5]), .B(rw), .Z(n6_adj_298)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3620_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_338 (.A(read_value[5]), .B(read_value_adj_186[5]), 
         .C(n52), .D(n64), .Z(n10_adj_300)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_338.init = 16'heca0;
    LUT4 i1_2_lut (.A(\register_addr[4] ), .B(\register_addr[5] ), .Z(n30427)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_339 (.A(\read_value[21]_adj_150 ), .B(read_value[21]), 
         .C(n32375), .D(n52), .Z(n8_adj_291)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_339.init = 16'heca0;
    PFUMX i25184 (.BLUT(n32220), .ALUT(n32219), .C0(\register_addr[1] ), 
          .Z(n32221));
    L6MUX21 i25178 (.D0(n32190), .D1(n32187), .SD(\register_addr[2] ), 
            .Z(n32191));
    PFUMX i24916 (.BLUT(n31486), .ALUT(n31485), .C0(\register_addr[1] ), 
          .Z(n31487));
    L6MUX21 i24938 (.D0(n31521), .D1(n31518), .SD(\register_addr[2] ), 
            .Z(n31522));
    PFUMX i25176 (.BLUT(n32189), .ALUT(n32188), .C0(\register_addr[1] ), 
          .Z(n32190));
    PFUMX i24936 (.BLUT(n31520), .ALUT(n31519), .C0(\register_addr[1] ), 
          .Z(n31521));
    PFUMX i25173 (.BLUT(n32186), .ALUT(n32185), .C0(\register_addr[1] ), 
          .Z(n32187));
    LUT4 i5_4_lut_adj_340 (.A(databus_out[20]), .B(n10_adj_307), .C(n2_adj_151), 
         .D(rw), .Z(databus[20])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_340.init = 16'hfcfe;
    LUT4 i1_4_lut (.A(\select[2] ), .B(read_size_c[0]), .C(\read_size[0]_adj_152 ), 
         .D(\select[7] ), .Z(n5)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i2_4_lut_adj_341 (.A(read_size[0]), .B(n25), .C(\select[1] ), 
         .D(n32439), .Z(n6_adj_153)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_341.init = 16'heca0;
    LUT4 i5_4_lut_adj_342 (.A(databus_out[31]), .B(n10_adj_312), .C(n2_adj_154), 
         .D(rw), .Z(databus[31])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_342.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_343 (.A(\read_value[31]_adj_155 ), .B(n8_adj_314), 
         .C(n1_adj_156), .D(n32472), .Z(n10_adj_312)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_343.init = 16'hfefc;
    LUT4 i2_4_lut_adj_344 (.A(\read_value[31]_adj_157 ), .B(read_value[31]), 
         .C(n32375), .D(n52), .Z(n8_adj_314)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_344.init = 16'heca0;
    LUT4 i1_4_lut_adj_345 (.A(read_size[2]), .B(n24), .C(\select[1] ), 
         .D(n32439), .Z(\reg_size[2] )) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_345.init = 16'heca0;
    LUT4 i5_4_lut_adj_346 (.A(databus_out[28]), .B(n10_adj_319), .C(n2_adj_158), 
         .D(rw), .Z(databus[28])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_346.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_347 (.A(\read_value[28]_adj_159 ), .B(n8_adj_321), 
         .C(n1_adj_160), .D(n32472), .Z(n10_adj_319)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_347.init = 16'hfefc;
    LUT4 i2_4_lut_adj_348 (.A(\read_value[28]_adj_161 ), .B(read_value[28]), 
         .C(n32375), .D(n52), .Z(n8_adj_321)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_348.init = 16'heca0;
    L6MUX21 i25150 (.D0(n32107), .D1(n32104), .SD(\register_addr[2] ), 
            .Z(n32108));
    PFUMX i25148 (.BLUT(n32106), .ALUT(n32105), .C0(\register_addr[1] ), 
          .Z(n32107));
    LUT4 i1_2_lut_adj_349 (.A(\register_addr[0] ), .B(\register_addr[1] ), 
         .Z(n30401)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_349.init = 16'h8888;
    LUT4 i4_4_lut_adj_350 (.A(\read_value[20]_adj_162 ), .B(n8_adj_325), 
         .C(n1_adj_163), .D(n32472), .Z(n10_adj_307)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_350.init = 16'hfefc;
    PFUMX i25145 (.BLUT(n32103), .ALUT(n32102), .C0(\register_addr[1] ), 
          .Z(n32104));
    LUT4 i7_4_lut_adj_351 (.A(n13_adj_327), .B(n4_adj_164), .C(n12_adj_329), 
         .D(n6_adj_330), .Z(databus[4])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_351.init = 16'hfffe;
    LUT4 i5_4_lut_adj_352 (.A(\read_value[4]_adj_165 ), .B(n10_adj_332), 
         .C(n7_adj_163), .D(n32374), .Z(n13_adj_327)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_352.init = 16'hfefc;
    LUT4 i4_4_lut_adj_353 (.A(\read_value[4]_adj_166 ), .B(\read_value[4]_adj_167 ), 
         .C(n32376), .D(n32472), .Z(n12_adj_329)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_353.init = 16'heca0;
    LUT4 Select_3621_i6_2_lut (.A(databus_out[4]), .B(rw), .Z(n6_adj_330)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3621_i6_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_354 (.A(read_value[4]), .B(read_value_adj_186[4]), 
         .C(n52), .D(n64), .Z(n10_adj_332)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_354.init = 16'heca0;
    PFUMX i24933 (.BLUT(n31517), .ALUT(n31516), .C0(\register_addr[1] ), 
          .Z(n31518));
    LUT4 i2_4_lut_adj_355 (.A(\read_value[20]_adj_168 ), .B(read_value[20]), 
         .C(n32375), .D(n52), .Z(n8_adj_325)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_355.init = 16'heca0;
    LUT4 i5_4_lut_adj_356 (.A(databus_out[27]), .B(n10_adj_339), .C(n2_adj_169), 
         .D(rw), .Z(databus[27])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_356.init = 16'hfcfe;
    L6MUX21 i25105 (.D0(n31902), .D1(n31899), .SD(\register_addr[2] ), 
            .Z(n31903));
    L6MUX21 i24921 (.D0(n31490), .D1(n31487), .SD(\register_addr[2] ), 
            .Z(n31491));
    LUT4 i4_4_lut_adj_357 (.A(\read_value[27]_adj_170 ), .B(n8_adj_341), 
         .C(n1_adj_171), .D(n32472), .Z(n10_adj_339)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_357.init = 16'hfefc;
    LUT4 i2_4_lut_adj_358 (.A(\read_value[27]_adj_172 ), .B(read_value[27]), 
         .C(n32375), .D(n52), .Z(n8_adj_341)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_358.init = 16'heca0;
    PFUMX i25101 (.BLUT(n31898), .ALUT(n31897), .C0(\register_addr[1] ), 
          .Z(n31899));
    LUT4 i5_4_lut_adj_359 (.A(databus_out[26]), .B(n10_adj_345), .C(n2_adj_173), 
         .D(rw), .Z(databus[26])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_359.init = 16'hfcfe;
    LUT4 i4_4_lut_adj_360 (.A(\read_value[26]_adj_174 ), .B(n8_adj_347), 
         .C(n1_adj_175), .D(n32472), .Z(n10_adj_345)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_360.init = 16'hfefc;
    PFUMX i25103 (.BLUT(n31901), .ALUT(n31900), .C0(\register_addr[1] ), 
          .Z(n31902));
    LUT4 i2_4_lut_adj_361 (.A(\read_value[26]_adj_176 ), .B(read_value[26]), 
         .C(n32375), .D(n52), .Z(n8_adj_347)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_361.init = 16'heca0;
    LUT4 i7_4_lut_adj_362 (.A(n13_adj_351), .B(n4_adj_177), .C(n12_adj_353), 
         .D(n6_adj_354), .Z(databus[3])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_362.init = 16'hfffe;
    LUT4 i5_4_lut_adj_363 (.A(\read_value[3]_adj_178 ), .B(n10_adj_356), 
         .C(n7_adj_162), .D(n32374), .Z(n13_adj_351)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_363.init = 16'hfefc;
    LUT4 i4_4_lut_adj_364 (.A(\read_value[3]_adj_179 ), .B(\read_value[3]_adj_180 ), 
         .C(n32376), .D(n32472), .Z(n12_adj_353)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_364.init = 16'heca0;
    LUT4 Select_3622_i6_2_lut (.A(databus_out[3]), .B(rw), .Z(n6_adj_354)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3622_i6_2_lut.init = 16'h2222;
    LUT4 i5_4_lut_adj_365 (.A(databus_out[25]), .B(n10_adj_359), .C(n2_adj_181), 
         .D(rw), .Z(databus[25])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_365.init = 16'hfcfe;
    LUT4 i2_4_lut_adj_366 (.A(read_value[3]), .B(read_value_adj_186[3]), 
         .C(n52), .D(n64), .Z(n10_adj_356)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_366.init = 16'heca0;
    LUT4 i4_4_lut_adj_367 (.A(\read_value[25]_adj_182 ), .B(n8_adj_363), 
         .C(n1_adj_183), .D(n32472), .Z(n10_adj_359)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_367.init = 16'hfefc;
    LUT4 i2_4_lut_adj_368 (.A(\read_value[25]_adj_184 ), .B(read_value[25]), 
         .C(n32375), .D(n52), .Z(n8_adj_363)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_368.init = 16'heca0;
    PFUMX i24919 (.BLUT(n31489), .ALUT(n31488), .C0(\register_addr[1] ), 
          .Z(n31490));
    PWMReceiver recv_ch8 (.n1054(n1054), .debug_c_c(debug_c_c), .n28324(n28324), 
            .GND_net(GND_net), .n32341(n32341), .rc_ch8_c(rc_ch8_c), .n31024(n31024), 
            .n30913(n30913), .\register[6] ({\register[6] }), .n12030(n12030)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(259[14] 263[36])
    PWMReceiver_U1 recv_ch7 (.n31005(n31005), .n1039(n1039), .debug_c_c(debug_c_c), 
            .n28308(n28308), .GND_net(GND_net), .n32341(n32341), .rc_ch7_c(rc_ch7_c), 
            .n30995(n30995), .\register[5] ({\register[5] }), .n12031(n12031)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(254[14] 258[36])
    PWMReceiver_U2 recv_ch4 (.\register[4] ({\register[4] }), .debug_c_c(debug_c_c), 
            .n32341(n32341), .GND_net(GND_net), .n30929(n30929), .rc_ch4_c(rc_ch4_c), 
            .n1024(n1024), .n28304(n28304)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(249[14] 253[36])
    PWMReceiver_U3 recv_ch3 (.debug_c_c(debug_c_c), .n32341(n32341), .GND_net(GND_net), 
            .\register[3] ({\register[3] }), .n12138(n12138), .n31000(n31000), 
            .n30969(n30969), .n1009(n1009), .n28317(n28317), .rc_ch3_c(rc_ch3_c)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(244[14] 248[36])
    PWMReceiver_U4 recv_ch2 (.n1000(n1000), .n988(n988), .n32341(n32341), 
            .debug_c_c(debug_c_c), .GND_net(GND_net), .\register[2] ({\register[2] }), 
            .n32336(n32336), .n14446(n14446), .n994(n994), .rc_ch2_c(rc_ch2_c), 
            .n54(n54), .n4(n4_adj_185)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(239[14] 243[36])
    PWMReceiver_U5 recv_ch1 (.debug_c_c(debug_c_c), .n32341(n32341), .GND_net(GND_net), 
            .\register[1] ({\register[1] }), .n12841(n12841), .n31049(n31049), 
            .n979(n979), .n28312(n28312), .rc_ch1_c(rc_ch1_c), .n30911(n30911)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(234[17] 238[36])
    
endmodule
//
// Verilog Description of module PWMReceiver
//

module PWMReceiver (n1054, debug_c_c, n28324, GND_net, n32341, rc_ch8_c, 
            n31024, n30913, \register[6] , n12030) /* synthesis syn_module_defined=1 */ ;
    output n1054;
    input debug_c_c;
    input n28324;
    input GND_net;
    input n32341;
    input rc_ch8_c;
    output n31024;
    output n30913;
    output [7:0]\register[6] ;
    input n12030;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    
    wire n11840, n4, n28401, n32456, n4_adj_133, n1060, n1048, 
        n30459, n32391, n30431, n28171, n10, n30656, n32393, n30493, 
        n32367, n30506;
    wire [7:0]n943;
    
    wire n30097;
    wire [7:0]n43;
    
    wire n32509, n32457, n32508, n28482, n32507, n32510, n32419, 
        n32441, n28353, n32420, n32506, n28321, n30148, n54, n32459, 
        n4_adj_134, n20244, n6, n32458, n30505;
    wire [15:0]n116;
    
    wire n14198, n14, n24, n27321, n27320, n27319, n27318, n27317, 
        n27316, n27315, n27314, n27609, n27608, n27607, n27606;
    
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n11840), .D(n4), 
         .Z(n28401)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_4_lut (.A(count[5]), .B(count[9]), .C(n32456), .D(n4_adj_133), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hfcec;
    LUT4 i1_2_lut (.A(n1060), .B(n1048), .Z(n30459)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n32391), .C(n30431), 
         .D(n28171), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i24299_3_lut_4_lut (.A(count[8]), .B(n32391), .C(n28171), .D(n30431), 
         .Z(n30656)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i24299_3_lut_4_lut.init = 16'hfeee;
    LUT4 i24771_3_lut_4_lut_4_lut (.A(n32393), .B(n30493), .C(n32367), 
         .D(n28171), .Z(n30506)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i24771_3_lut_4_lut_4_lut.init = 16'h1110;
    LUT4 i14246_2_lut (.A(n943[0]), .B(n30097), .Z(n43[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14246_2_lut.init = 16'h2222;
    LUT4 i3_3_lut_4_lut (.A(count[8]), .B(n32509), .C(n32457), .D(n32508), 
         .Z(n28482)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32508), .B(n32509), .C(n32507), .D(count[0]), 
         .Z(n30431)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_325_3_lut_4_lut (.A(n32510), .B(count[13]), .C(n11840), 
         .D(count[12]), .Z(n32419)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_325_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_273_3_lut_4_lut (.A(n11840), .B(n32441), .C(count[8]), 
         .D(count[9]), .Z(n32367)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_273_3_lut_4_lut.init = 16'hfffe;
    LUT4 i14730_2_lut_rep_326 (.A(n28353), .B(count[9]), .Z(n32420)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14730_2_lut_rep_326.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_257 (.A(n28353), .B(count[9]), .C(n32441), 
         .D(n11840), .Z(n30493)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_257.init = 16'hfff8;
    FD1P3IX valid_48 (.D(n30506), .SP(n28324), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1054));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch8_c), .SP(n32341), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1060));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1060), .SP(n32341), .CK(debug_c_c), .Q(n1048));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i24756_4_lut (.A(n32510), .B(n32506), .C(n28401), .D(n28321), 
         .Z(n31024)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i24756_4_lut.init = 16'h3233;
    LUT4 i1_4_lut_adj_258 (.A(n30656), .B(n30459), .C(n11840), .D(n30148), 
         .Z(n28321)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_258.init = 16'hcecc;
    LUT4 i3_4_lut (.A(n54), .B(n32420), .C(n30097), .D(n32441), .Z(n30148)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_adj_259 (.A(count[11]), .B(count[10]), .Z(n11840)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_259.init = 16'heeee;
    LUT4 i1_2_lut_rep_297_3_lut_4_lut (.A(count[12]), .B(n32459), .C(count[9]), 
         .D(n11840), .Z(n32391)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_297_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_260 (.A(count[4]), .B(count[5]), .C(n4_adj_134), 
         .D(n32509), .Z(n28171)) /* synthesis lut_function=(A (B (D))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i2_4_lut_adj_260.init = 16'hc800;
    LUT4 i3_4_lut_adj_261 (.A(count[7]), .B(count[8]), .C(n20244), .D(count[6]), 
         .Z(n28353)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_261.init = 16'hfffe;
    LUT4 i14512_4_lut (.A(count[0]), .B(n32508), .C(n6), .D(count[3]), 
         .Z(n20244)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i14512_4_lut.init = 16'hccc8;
    LUT4 i2_2_lut (.A(count[1]), .B(count[2]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_262 (.A(n32391), .B(count[8]), .C(n32507), .D(n32458), 
         .Z(n30097)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i1_4_lut_adj_262.init = 16'hfbbb;
    LUT4 n28482_bdd_4_lut (.A(n28482), .B(count[9]), .C(n28353), .D(n32419), 
         .Z(n54)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A ((C+(D))+!B))) */ ;
    defparam n28482_bdd_4_lut.init = 16'h002e;
    LUT4 i5_2_lut_rep_412 (.A(n1048), .B(n1060), .Z(n32506)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i5_2_lut_rep_412.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_263 (.A(n1048), .B(n1060), .C(n28401), 
         .D(n32510), .Z(n30505)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i1_2_lut_3_lut_4_lut_adj_263.init = 16'hfff4;
    LUT4 i2_3_lut_rep_413 (.A(count[2]), .B(count[3]), .C(count[1]), .Z(n32507)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_rep_413.init = 16'h8080;
    LUT4 i1_2_lut_rep_363_4_lut (.A(count[2]), .B(count[3]), .C(count[1]), 
         .D(count[0]), .Z(n32457)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_363_4_lut.init = 16'h8000;
    LUT4 i14028_2_lut_rep_414 (.A(count[5]), .B(count[4]), .Z(n32508)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14028_2_lut_rep_414.init = 16'h8888;
    LUT4 i1_2_lut_rep_415 (.A(count[6]), .B(count[7]), .Z(n32509)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_415.init = 16'h8888;
    LUT4 i1_2_lut_rep_362_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n32456)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_362_3_lut.init = 16'h8080;
    LUT4 i2_2_lut_rep_364_3_lut_4_lut (.A(count[6]), .B(count[7]), .C(count[4]), 
         .D(count[5]), .Z(n32458)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_2_lut_rep_364_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut (.A(count[1]), .B(count[2]), .C(count[3]), .Z(n4_adj_134)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[1]), .B(count[2]), .C(count[3]), .D(count[4]), 
         .Z(n4_adj_133)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff80;
    LUT4 i1_2_lut_rep_416 (.A(count[15]), .B(count[14]), .Z(n32510)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_416.init = 16'heeee;
    LUT4 i2_2_lut_rep_347_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(count[12]), 
         .D(count[13]), .Z(n32441)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_2_lut_rep_347_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_299_3_lut (.A(count[15]), .B(count[14]), .C(n28401), 
         .Z(n32393)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_299_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_365_3_lut (.A(count[15]), .B(count[14]), .C(count[13]), 
         .Z(n32459)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_365_3_lut.init = 16'hfefe;
    LUT4 i24645_4_lut (.A(n54), .B(n30459), .C(n30097), .D(n10), .Z(n30913)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i24645_4_lut.init = 16'h3323;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    LUT4 i7_4_lut (.A(n1048), .B(n14), .C(n32459), .D(n1060), .Z(n14198)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i7_4_lut.init = 16'h0008;
    LUT4 i6_4_lut (.A(count[12]), .B(n24), .C(n11840), .D(n32341), .Z(n14)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i6_4_lut.init = 16'h0400;
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    LUT4 i31_3_lut (.A(n28482), .B(n28353), .C(count[9]), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i31_3_lut.init = 16'h3a3a;
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    LUT4 i14444_2_lut (.A(n943[1]), .B(n30097), .Z(n43[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14444_2_lut.init = 16'h2222;
    LUT4 i14445_2_lut (.A(n943[2]), .B(n30097), .Z(n43[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14445_2_lut.init = 16'h2222;
    LUT4 i14446_2_lut (.A(n943[3]), .B(n30097), .Z(n43[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14446_2_lut.init = 16'h2222;
    LUT4 i14447_2_lut (.A(n943[4]), .B(n30097), .Z(n43[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14447_2_lut.init = 16'h2222;
    LUT4 i14448_2_lut (.A(n943[5]), .B(n30097), .Z(n43[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14448_2_lut.init = 16'h2222;
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n12030), .PD(n14198), .CK(debug_c_c), 
            .Q(\register[6] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i14449_2_lut (.A(n943[6]), .B(n30097), .Z(n43[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14449_2_lut.init = 16'h2222;
    LUT4 i14450_2_lut (.A(n943[7]), .B(n30097), .Z(n43[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14450_2_lut.init = 16'h2222;
    CCU2D add_1493_17 (.A0(count[15]), .B0(n32506), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27321), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_17.INIT0 = 16'hd222;
    defparam add_1493_17.INIT1 = 16'h0000;
    defparam add_1493_17.INJECT1_0 = "NO";
    defparam add_1493_17.INJECT1_1 = "NO";
    CCU2D add_1493_15 (.A0(count[13]), .B0(n32506), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n32506), .C1(GND_net), .D1(GND_net), .CIN(n27320), 
          .COUT(n27321), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_15.INIT0 = 16'hd222;
    defparam add_1493_15.INIT1 = 16'hd222;
    defparam add_1493_15.INJECT1_0 = "NO";
    defparam add_1493_15.INJECT1_1 = "NO";
    CCU2D add_1493_13 (.A0(count[11]), .B0(n32506), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n32506), .C1(GND_net), .D1(GND_net), .CIN(n27319), 
          .COUT(n27320), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_13.INIT0 = 16'hd222;
    defparam add_1493_13.INIT1 = 16'hd222;
    defparam add_1493_13.INJECT1_0 = "NO";
    defparam add_1493_13.INJECT1_1 = "NO";
    CCU2D add_1493_11 (.A0(count[9]), .B0(n32506), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n32506), .C1(GND_net), .D1(GND_net), .CIN(n27318), 
          .COUT(n27319), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_11.INIT0 = 16'hd222;
    defparam add_1493_11.INIT1 = 16'hd222;
    defparam add_1493_11.INJECT1_0 = "NO";
    defparam add_1493_11.INJECT1_1 = "NO";
    CCU2D add_1493_9 (.A0(count[7]), .B0(n32506), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n32506), .C1(GND_net), .D1(GND_net), .CIN(n27317), 
          .COUT(n27318), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_9.INIT0 = 16'hd222;
    defparam add_1493_9.INIT1 = 16'hd222;
    defparam add_1493_9.INJECT1_0 = "NO";
    defparam add_1493_9.INJECT1_1 = "NO";
    CCU2D add_1493_7 (.A0(count[5]), .B0(n32506), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n32506), .C1(GND_net), .D1(GND_net), .CIN(n27316), 
          .COUT(n27317), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_7.INIT0 = 16'hd222;
    defparam add_1493_7.INIT1 = 16'hd222;
    defparam add_1493_7.INJECT1_0 = "NO";
    defparam add_1493_7.INJECT1_1 = "NO";
    CCU2D add_1493_5 (.A0(count[3]), .B0(n32506), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n32506), .C1(GND_net), .D1(GND_net), .CIN(n27315), 
          .COUT(n27316), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_5.INIT0 = 16'hd222;
    defparam add_1493_5.INIT1 = 16'hd222;
    defparam add_1493_5.INJECT1_0 = "NO";
    defparam add_1493_5.INJECT1_1 = "NO";
    CCU2D add_1493_3 (.A0(count[1]), .B0(n32506), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n32506), .C1(GND_net), .D1(GND_net), .CIN(n27314), 
          .COUT(n27315), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_3.INIT0 = 16'hd222;
    defparam add_1493_3.INIT1 = 16'hd222;
    defparam add_1493_3.INJECT1_0 = "NO";
    defparam add_1493_3.INJECT1_1 = "NO";
    CCU2D add_1493_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n30505), .B1(n1060), .C1(count[0]), .D1(n1048), .COUT(n27314), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1493_1.INIT0 = 16'hF000;
    defparam add_1493_1.INIT1 = 16'ha565;
    defparam add_1493_1.INJECT1_0 = "NO";
    defparam add_1493_1.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27609), 
          .S0(n943[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_61_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_9.INIT1 = 16'h0000;
    defparam sub_61_add_2_9.INJECT1_0 = "NO";
    defparam sub_61_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27608), 
          .COUT(n27609), .S0(n943[5]), .S1(n943[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_61_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_61_add_2_7.INJECT1_0 = "NO";
    defparam sub_61_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27607), 
          .COUT(n27608), .S0(n943[3]), .S1(n943[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_61_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_61_add_2_5.INJECT1_0 = "NO";
    defparam sub_61_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27606), 
          .COUT(n27607), .S0(n943[1]), .S1(n943[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_61_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_61_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_61_add_2_3.INJECT1_0 = "NO";
    defparam sub_61_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_61_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27606), 
          .S1(n943[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_61_add_2_1.INIT0 = 16'hF000;
    defparam sub_61_add_2_1.INIT1 = 16'h5555;
    defparam sub_61_add_2_1.INJECT1_0 = "NO";
    defparam sub_61_add_2_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMReceiver_U1
//

module PWMReceiver_U1 (n31005, n1039, debug_c_c, n28308, GND_net, 
            n32341, rc_ch7_c, n30995, \register[5] , n12031) /* synthesis syn_module_defined=1 */ ;
    output n31005;
    output n1039;
    input debug_c_c;
    input n28308;
    input GND_net;
    input n32341;
    input rc_ch7_c;
    output n30995;
    output [7:0]\register[5] ;
    input n12031;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n32501, n32499, n28466, n28307, n32436, n30480, n12, 
        n8, n32415, n30565, n32414, n4, n54, n30111;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    
    wire n6, n11927, n1045, n1033, n32500, n32437, n28374, n6_adj_131, 
        n28245, n4_adj_132;
    wire [7:0]n934;
    wire [7:0]n43;
    
    wire n32502, n28188, n32438, n32453, n30491, n30451, n29791, 
        n30490, n32388, n10, n30160, n14177, n30671, n24;
    wire [15:0]n116;
    
    wire n27329, n27328, n27327, n27326, n27325, n27324, n27323, 
        n27322, n27613, n27612, n27611, n27610;
    
    LUT4 i24737_4_lut (.A(n32501), .B(n32499), .C(n28466), .D(n28307), 
         .Z(n31005)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i24737_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n32436), .B(n30480), .C(n12), .D(n8), .Z(n28307)) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hdccc;
    LUT4 i5_4_lut (.A(n32415), .B(n30565), .C(n32414), .D(n4), .Z(n12)) /* synthesis lut_function=(!(A (B)+!A (B+!(C (D))))) */ ;
    defparam i5_4_lut.init = 16'h3222;
    LUT4 i1_2_lut (.A(n54), .B(n30111), .Z(n8)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i1_4_lut_adj_240 (.A(count[4]), .B(count[5]), .C(count[3]), .D(n6), 
         .Z(n4)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_240.init = 16'hccc8;
    LUT4 i2_2_lut (.A(count[1]), .B(count[2]), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i24213_4_lut (.A(count[12]), .B(n11927), .C(n32501), .D(count[13]), 
         .Z(n30565)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24213_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_241 (.A(count[11]), .B(count[10]), .Z(n11927)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_adj_241.init = 16'heeee;
    LUT4 i1_2_lut_adj_242 (.A(n1045), .B(n1033), .Z(n30480)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_242.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_343_4_lut (.A(count[3]), .B(n6), .C(n32500), .D(count[0]), 
         .Z(n32437)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_343_4_lut.init = 16'h8000;
    LUT4 i3_4_lut (.A(n28374), .B(n6_adj_131), .C(count[8]), .D(n32500), 
         .Z(n28245)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i3_4_lut.init = 16'hfefc;
    LUT4 i3_4_lut_adj_243 (.A(count[0]), .B(count[1]), .C(count[3]), .D(count[2]), 
         .Z(n28374)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_243.init = 16'hfffe;
    LUT4 i2_2_lut_adj_244 (.A(count[6]), .B(count[7]), .Z(n6_adj_131)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_2_lut_adj_244.init = 16'heeee;
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n11927), .D(n4_adj_132), 
         .Z(n28466)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_2_lut_adj_245 (.A(n30111), .B(n934[5]), .Z(n43[5])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_245.init = 16'h4444;
    LUT4 i1_4_lut_adj_246 (.A(n32502), .B(count[9]), .C(n28188), .D(count[8]), 
         .Z(n4_adj_132)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_246.init = 16'heccc;
    LUT4 i1_2_lut_adj_247 (.A(n30111), .B(n934[6]), .Z(n43[6])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_247.init = 16'h4444;
    LUT4 i1_2_lut_adj_248 (.A(n30111), .B(n934[7]), .Z(n43[7])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_248.init = 16'h4444;
    LUT4 i2_4_lut_adj_249 (.A(count[5]), .B(count[4]), .C(n6), .D(count[3]), 
         .Z(n28188)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_249.init = 16'hfeee;
    LUT4 i1_4_lut_adj_250 (.A(n32438), .B(count[8]), .C(n32502), .D(n32453), 
         .Z(n30111)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i1_4_lut_adj_250.init = 16'hfbbb;
    FD1P3IX valid_48 (.D(n30491), .SP(n28308), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1039));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch7_c), .SP(n32341), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1045));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n1045), .SP(n32341), .CK(debug_c_c), .Q(n1033));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i14571_2_lut_rep_342 (.A(n28245), .B(count[9]), .Z(n32436)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14571_2_lut_rep_342.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(n28245), .B(count[9]), .C(n30565), .Z(n30451)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[0]), .B(n32453), .C(n32502), .D(count[8]), 
         .Z(n29791)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h8000;
    LUT4 n29791_bdd_4_lut_25308 (.A(n29791), .B(count[9]), .C(n28245), 
         .D(n30565), .Z(n54)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A ((C+(D))+!B))) */ ;
    defparam n29791_bdd_4_lut_25308.init = 16'h002e;
    LUT4 i1_2_lut_rep_344 (.A(count[9]), .B(n30565), .Z(n32438)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_344.init = 16'heeee;
    LUT4 i1_2_lut_rep_321_3_lut (.A(count[9]), .B(n30565), .C(count[8]), 
         .Z(n32415)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_321_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_adj_251 (.A(n30111), .B(n934[2]), .Z(n43[2])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_251.init = 16'h4444;
    LUT4 i5_2_lut_rep_405 (.A(n1033), .B(n1045), .Z(n32499)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i5_2_lut_rep_405.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n1033), .B(n1045), .C(n28466), .D(n32501), 
         .Z(n30490)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff4;
    LUT4 i1_2_lut_rep_406 (.A(count[4]), .B(count[5]), .Z(n32500)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_406.init = 16'h8888;
    LUT4 i3_3_lut_rep_359_4_lut (.A(count[4]), .B(count[5]), .C(n6), .D(count[3]), 
         .Z(n32453)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_3_lut_rep_359_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_407 (.A(count[15]), .B(count[14]), .Z(n32501)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_407.init = 16'heeee;
    LUT4 i1_2_lut_rep_408 (.A(count[6]), .B(count[7]), .Z(n32502)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_408.init = 16'h8888;
    LUT4 i1_2_lut_rep_320_3_lut_4_lut (.A(count[6]), .B(count[7]), .C(n32453), 
         .D(count[0]), .Z(n32414)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_320_3_lut_4_lut.init = 16'h8000;
    LUT4 i24769_3_lut_3_lut_4_lut (.A(n32501), .B(n28466), .C(n32388), 
         .D(n30451), .Z(n30491)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i24769_3_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i24727_4_lut (.A(n54), .B(n30480), .C(n30111), .D(n10), .Z(n30995)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i24727_4_lut.init = 16'h3323;
    LUT4 i3_4_lut_adj_252 (.A(n32501), .B(n30160), .C(n11927), .D(n32341), 
         .Z(n14177)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut_adj_252.init = 16'h0400;
    LUT4 i1_2_lut_adj_253 (.A(n30111), .B(n934[3]), .Z(n43[3])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_253.init = 16'h4444;
    LUT4 i4_4_lut (.A(n30671), .B(n24), .C(n1033), .D(n1045), .Z(n30160)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i4_4_lut.init = 16'h0040;
    LUT4 i24313_2_lut (.A(count[13]), .B(count[12]), .Z(n30671)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24313_2_lut.init = 16'heeee;
    LUT4 i31_3_lut (.A(n29791), .B(n28245), .C(count[9]), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i31_3_lut.init = 16'h3a3a;
    LUT4 i1_2_lut_adj_254 (.A(n30111), .B(n934[0]), .Z(n43[0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_254.init = 16'h4444;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_255 (.A(n30111), .B(n934[4]), .Z(n43[4])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_255.init = 16'h4444;
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n12031), .PD(n14177), .CK(debug_c_c), 
            .Q(\register[5] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    CCU2D add_1489_17 (.A0(count[15]), .B0(n32499), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27329), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_17.INIT0 = 16'hd222;
    defparam add_1489_17.INIT1 = 16'h0000;
    defparam add_1489_17.INJECT1_0 = "NO";
    defparam add_1489_17.INJECT1_1 = "NO";
    CCU2D add_1489_15 (.A0(count[13]), .B0(n32499), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n32499), .C1(GND_net), .D1(GND_net), .CIN(n27328), 
          .COUT(n27329), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_15.INIT0 = 16'hd222;
    defparam add_1489_15.INIT1 = 16'hd222;
    defparam add_1489_15.INJECT1_0 = "NO";
    defparam add_1489_15.INJECT1_1 = "NO";
    CCU2D add_1489_13 (.A0(count[11]), .B0(n32499), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n32499), .C1(GND_net), .D1(GND_net), .CIN(n27327), 
          .COUT(n27328), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_13.INIT0 = 16'hd222;
    defparam add_1489_13.INIT1 = 16'hd222;
    defparam add_1489_13.INJECT1_0 = "NO";
    defparam add_1489_13.INJECT1_1 = "NO";
    CCU2D add_1489_11 (.A0(count[9]), .B0(n32499), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n32499), .C1(GND_net), .D1(GND_net), .CIN(n27326), 
          .COUT(n27327), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_11.INIT0 = 16'hd222;
    defparam add_1489_11.INIT1 = 16'hd222;
    defparam add_1489_11.INJECT1_0 = "NO";
    defparam add_1489_11.INJECT1_1 = "NO";
    CCU2D add_1489_9 (.A0(count[7]), .B0(n32499), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n32499), .C1(GND_net), .D1(GND_net), .CIN(n27325), 
          .COUT(n27326), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_9.INIT0 = 16'hd222;
    defparam add_1489_9.INIT1 = 16'hd222;
    defparam add_1489_9.INJECT1_0 = "NO";
    defparam add_1489_9.INJECT1_1 = "NO";
    CCU2D add_1489_7 (.A0(count[5]), .B0(n32499), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n32499), .C1(GND_net), .D1(GND_net), .CIN(n27324), 
          .COUT(n27325), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_7.INIT0 = 16'hd222;
    defparam add_1489_7.INIT1 = 16'hd222;
    defparam add_1489_7.INJECT1_0 = "NO";
    defparam add_1489_7.INJECT1_1 = "NO";
    CCU2D add_1489_5 (.A0(count[3]), .B0(n32499), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n32499), .C1(GND_net), .D1(GND_net), .CIN(n27323), 
          .COUT(n27324), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_5.INIT0 = 16'hd222;
    defparam add_1489_5.INIT1 = 16'hd222;
    defparam add_1489_5.INJECT1_0 = "NO";
    defparam add_1489_5.INJECT1_1 = "NO";
    CCU2D add_1489_3 (.A0(count[1]), .B0(n32499), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n32499), .C1(GND_net), .D1(GND_net), .CIN(n27322), 
          .COUT(n27323), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_3.INIT0 = 16'hd222;
    defparam add_1489_3.INIT1 = 16'hd222;
    defparam add_1489_3.INJECT1_0 = "NO";
    defparam add_1489_3.INJECT1_1 = "NO";
    CCU2D add_1489_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n30490), .B1(n1045), .C1(count[0]), .D1(n1033), .COUT(n27322), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1489_1.INIT0 = 16'hF000;
    defparam add_1489_1.INIT1 = 16'ha565;
    defparam add_1489_1.INJECT1_0 = "NO";
    defparam add_1489_1.INJECT1_1 = "NO";
    CCU2D sub_60_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27613), 
          .S0(n934[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_60_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_9.INIT1 = 16'h0000;
    defparam sub_60_add_2_9.INJECT1_0 = "NO";
    defparam sub_60_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_60_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27612), 
          .COUT(n27613), .S0(n934[5]), .S1(n934[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_60_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_60_add_2_7.INJECT1_0 = "NO";
    defparam sub_60_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_60_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27611), 
          .COUT(n27612), .S0(n934[3]), .S1(n934[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_60_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_60_add_2_5.INJECT1_0 = "NO";
    defparam sub_60_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_60_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27610), 
          .COUT(n27611), .S0(n934[1]), .S1(n934[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_60_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_60_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_60_add_2_3.INJECT1_0 = "NO";
    defparam sub_60_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_60_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27610), 
          .S1(n934[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_60_add_2_1.INIT0 = 16'hF000;
    defparam sub_60_add_2_1.INIT1 = 16'h5555;
    defparam sub_60_add_2_1.INJECT1_0 = "NO";
    defparam sub_60_add_2_1.INJECT1_1 = "NO";
    LUT4 i10_3_lut_4_lut_4_lut (.A(n32502), .B(n32437), .C(n4), .D(n32415), 
         .Z(n10)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i10_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 i1_3_lut_rep_294_4_lut (.A(count[8]), .B(n32438), .C(n4), .D(n32502), 
         .Z(n32388)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_3_lut_rep_294_4_lut.init = 16'hfeee;
    LUT4 i1_2_lut_adj_256 (.A(n30111), .B(n934[1]), .Z(n43[1])) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_adj_256.init = 16'h4444;
    
endmodule
//
// Verilog Description of module PWMReceiver_U2
//

module PWMReceiver_U2 (\register[4] , debug_c_c, n32341, GND_net, n30929, 
            rc_ch4_c, n1024, n28304) /* synthesis syn_module_defined=1 */ ;
    output [7:0]\register[4] ;
    input debug_c_c;
    input n32341;
    input GND_net;
    output n30929;
    input rc_ch4_c;
    output n1024;
    input n28304;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n11987, n14143;
    wire [7:0]n43;
    
    wire n1018, n30158, n30573;
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    wire [15:0]n116;
    
    wire n32351, n28359, n1030, n30563, n32370, n30440, n32467, 
        n32397, n32466, n32396, n30414, n30500, n30499, n32446, 
        n4, n6, n32344, n32382, n32372, n20316, n30718, n11779, 
        n32430, n30465, n28378, n30467, n128_adj_129, n5, n6_adj_130, 
        n28375;
    wire [7:0]n925;
    
    wire n27337, n11813, n27336, n27335, n27334, n27333, n27332, 
        n27331, n27330, n27617, n27616, n27615, n27614;
    
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    LUT4 i3_4_lut (.A(n1018), .B(n32341), .C(n30158), .D(n30573), .Z(n14143)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut.init = 16'h0080;
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(n32351), .B(n28359), .C(count[9]), .D(n1030), 
         .Z(n30158)) /* synthesis lut_function=(!(A ((D)+!B)+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i2_4_lut.init = 16'h00c8;
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    LUT4 i2_2_lut_rep_276 (.A(count[0]), .B(n30563), .Z(n32370)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_rep_276.init = 16'h8888;
    LUT4 i24661_4_lut (.A(n30440), .B(n32467), .C(n32397), .D(n32466), 
         .Z(n30929)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i24661_4_lut.init = 16'h3031;
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_257_3_lut (.A(count[0]), .B(n30563), .C(count[8]), 
         .Z(n32351)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_257_3_lut.init = 16'h8080;
    LUT4 i24763_3_lut_4_lut_4_lut (.A(n32397), .B(n30573), .C(n32396), 
         .D(n30414), .Z(n30500)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i24763_3_lut_4_lut_4_lut.init = 16'h1110;
    LUT4 i1_2_lut_rep_372 (.A(n1030), .B(n1018), .Z(n32466)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_372.init = 16'hbbbb;
    LUT4 i24750_3_lut_3_lut_4_lut (.A(n1030), .B(n1018), .C(n28359), .D(n32341), 
         .Z(n11987)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i24750_3_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i5_2_lut_rep_373 (.A(n1018), .B(n1030), .Z(n32467)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i5_2_lut_rep_373.init = 16'h4444;
    LUT4 i1_2_lut_3_lut (.A(n1018), .B(n1030), .C(n32397), .Z(n30499)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i1_2_lut_3_lut.init = 16'hf4f4;
    LUT4 i1_2_lut_rep_352_3_lut (.A(count[6]), .B(count[7]), .C(count[5]), 
         .Z(n32446)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_rep_352_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_230 (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_3_lut_adj_230.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_4_lut (.A(count[6]), .B(count[7]), .C(count[2]), 
         .D(count[5]), .Z(n6)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1P3AX prev_in_46 (.D(n1030), .SP(n32341), .CK(debug_c_c), .Q(n1018));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch4_c), .SP(n32341), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1030));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_231 (.A(n32344), .B(n32382), .C(n32372), .D(n20316), 
         .Z(n28359)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i2_4_lut_adj_231.init = 16'heefe;
    LUT4 i3_4_lut_adj_232 (.A(n32396), .B(n30718), .C(n32370), .D(n30414), 
         .Z(n30440)) /* synthesis lut_function=(!(A (B)+!A (B+!(C (D))))) */ ;
    defparam i3_4_lut_adj_232.init = 16'h3222;
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_336 (.A(count[9]), .B(n11779), .Z(n32430)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_336.init = 16'heeee;
    LUT4 i1_3_lut_rep_288_4_lut (.A(count[9]), .B(n11779), .C(n30563), 
         .D(count[8]), .Z(n32382)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_3_lut_rep_288_4_lut.init = 16'h0100;
    LUT4 i2_4_lut_adj_233 (.A(n30465), .B(count[9]), .C(n28378), .D(n4), 
         .Z(n30467)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_233.init = 16'hfeee;
    LUT4 i2_4_lut_adj_234 (.A(count[3]), .B(count[4]), .C(n128_adj_129), 
         .D(count[5]), .Z(n28378)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_4_lut_adj_234.init = 16'hffec;
    LUT4 i1_2_lut_rep_302_3_lut (.A(count[9]), .B(n11779), .C(count[8]), 
         .Z(n32396)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_302_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut (.A(count[2]), .B(count[1]), .Z(n128_adj_129)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_278_3_lut_4_lut (.A(count[9]), .B(n11779), .C(n30414), 
         .D(count[8]), .Z(n32372)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_278_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21_3_lut_rep_250_4_lut (.A(count[8]), .B(n32370), .C(n32430), 
         .D(n30573), .Z(n32344)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i21_3_lut_rep_250_4_lut.init = 16'h00f8;
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    LUT4 i24219_4_lut (.A(n11779), .B(count[9]), .C(n5), .D(n6_adj_130), 
         .Z(n30573)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i24219_4_lut.init = 16'heeea;
    LUT4 i1_4_lut (.A(count[7]), .B(count[4]), .C(count[5]), .D(n28375), 
         .Z(n5)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_4_lut.init = 16'heaaa;
    LUT4 i2_2_lut (.A(count[8]), .B(count[6]), .Z(n6_adj_130)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_235 (.A(count[1]), .B(count[3]), .C(count[2]), .D(count[0]), 
         .Z(n28375)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i3_4_lut_adj_235.init = 16'hfffe;
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_236 (.A(n128_adj_129), .B(n32446), .C(count[4]), 
         .D(count[3]), .Z(n30414)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_4_lut_adj_236.init = 16'hccc8;
    LUT4 i14437_2_lut_4_lut (.A(count[8]), .B(n32430), .C(n30563), .D(n925[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14437_2_lut_4_lut.init = 16'h0200;
    LUT4 i14438_2_lut_4_lut (.A(count[8]), .B(n32430), .C(n30563), .D(n925[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14438_2_lut_4_lut.init = 16'h0200;
    FD1P3IX valid_48 (.D(n30500), .SP(n28304), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1024));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n11987), .PD(n14143), .CK(debug_c_c), 
            .Q(\register[4] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i14440_2_lut_4_lut (.A(count[8]), .B(n32430), .C(n30563), .D(n925[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14440_2_lut_4_lut.init = 16'h0200;
    LUT4 i24359_3_lut_4_lut (.A(n32351), .B(n30573), .C(n32430), .D(n32382), 
         .Z(n30718)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[13:39])
    defparam i24359_3_lut_4_lut.init = 16'hfffe;
    LUT4 i14577_2_lut_3_lut_4_lut (.A(count[8]), .B(n32430), .C(n30563), 
         .D(count[0]), .Z(n20316)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i14577_2_lut_3_lut_4_lut.init = 16'hfeee;
    CCU2D add_1485_17 (.A0(count[15]), .B0(n32467), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27337), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_17.INIT0 = 16'hd222;
    defparam add_1485_17.INIT1 = 16'h0000;
    defparam add_1485_17.INJECT1_0 = "NO";
    defparam add_1485_17.INJECT1_1 = "NO";
    LUT4 i1_4_lut_rep_303 (.A(n11813), .B(count[13]), .C(count[12]), .D(n30467), 
         .Z(n32397)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_rep_303.init = 16'heaaa;
    CCU2D add_1485_15 (.A0(count[13]), .B0(n32467), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n32467), .C1(GND_net), .D1(GND_net), .CIN(n27336), 
          .COUT(n27337), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_15.INIT0 = 16'hd222;
    defparam add_1485_15.INIT1 = 16'hd222;
    defparam add_1485_15.INJECT1_0 = "NO";
    defparam add_1485_15.INJECT1_1 = "NO";
    CCU2D add_1485_13 (.A0(count[11]), .B0(n32467), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n32467), .C1(GND_net), .D1(GND_net), .CIN(n27335), 
          .COUT(n27336), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_13.INIT0 = 16'hd222;
    defparam add_1485_13.INIT1 = 16'hd222;
    defparam add_1485_13.INJECT1_0 = "NO";
    defparam add_1485_13.INJECT1_1 = "NO";
    LUT4 i24211_4_lut (.A(count[1]), .B(count[3]), .C(n6), .D(count[4]), 
         .Z(n30563)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i24211_4_lut.init = 16'h8000;
    CCU2D add_1485_11 (.A0(count[9]), .B0(n32467), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n32467), .C1(GND_net), .D1(GND_net), .CIN(n27334), 
          .COUT(n27335), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_11.INIT0 = 16'hd222;
    defparam add_1485_11.INIT1 = 16'hd222;
    defparam add_1485_11.INJECT1_0 = "NO";
    defparam add_1485_11.INJECT1_1 = "NO";
    CCU2D add_1485_9 (.A0(count[7]), .B0(n32467), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n32467), .C1(GND_net), .D1(GND_net), .CIN(n27333), 
          .COUT(n27334), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_9.INIT0 = 16'hd222;
    defparam add_1485_9.INIT1 = 16'hd222;
    defparam add_1485_9.INJECT1_0 = "NO";
    defparam add_1485_9.INJECT1_1 = "NO";
    CCU2D add_1485_7 (.A0(count[5]), .B0(n32467), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n32467), .C1(GND_net), .D1(GND_net), .CIN(n27332), 
          .COUT(n27333), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_7.INIT0 = 16'hd222;
    defparam add_1485_7.INIT1 = 16'hd222;
    defparam add_1485_7.INJECT1_0 = "NO";
    defparam add_1485_7.INJECT1_1 = "NO";
    CCU2D add_1485_5 (.A0(count[3]), .B0(n32467), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n32467), .C1(GND_net), .D1(GND_net), .CIN(n27331), 
          .COUT(n27332), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_5.INIT0 = 16'hd222;
    defparam add_1485_5.INIT1 = 16'hd222;
    defparam add_1485_5.INJECT1_0 = "NO";
    defparam add_1485_5.INJECT1_1 = "NO";
    CCU2D add_1485_3 (.A0(count[1]), .B0(n32467), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n32467), .C1(GND_net), .D1(GND_net), .CIN(n27330), 
          .COUT(n27331), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_3.INIT0 = 16'hd222;
    defparam add_1485_3.INIT1 = 16'hd222;
    defparam add_1485_3.INJECT1_0 = "NO";
    defparam add_1485_3.INJECT1_1 = "NO";
    CCU2D add_1485_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n30499), .B1(n1030), .C1(count[0]), .D1(n1018), .COUT(n27330), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1485_1.INIT0 = 16'hF000;
    defparam add_1485_1.INIT1 = 16'ha565;
    defparam add_1485_1.INJECT1_0 = "NO";
    defparam add_1485_1.INJECT1_1 = "NO";
    LUT4 i3_4_lut_adj_237 (.A(count[12]), .B(count[13]), .C(n11813), .D(n30465), 
         .Z(n11779)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_237.init = 16'hfffe;
    LUT4 i14441_2_lut_4_lut (.A(count[8]), .B(n32430), .C(n30563), .D(n925[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14441_2_lut_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_adj_238 (.A(count[15]), .B(count[14]), .Z(n11813)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_238.init = 16'heeee;
    CCU2D sub_59_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27617), 
          .S0(n925[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_59_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_9.INIT1 = 16'h0000;
    defparam sub_59_add_2_9.INJECT1_0 = "NO";
    defparam sub_59_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_59_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27616), 
          .COUT(n27617), .S0(n925[5]), .S1(n925[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_59_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_59_add_2_7.INJECT1_0 = "NO";
    defparam sub_59_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_59_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27615), 
          .COUT(n27616), .S0(n925[3]), .S1(n925[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_59_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_59_add_2_5.INJECT1_0 = "NO";
    defparam sub_59_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_59_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27614), 
          .COUT(n27615), .S0(n925[1]), .S1(n925[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_59_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_59_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_59_add_2_3.INJECT1_0 = "NO";
    defparam sub_59_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_59_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27614), 
          .S1(n925[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_59_add_2_1.INIT0 = 16'hF000;
    defparam sub_59_add_2_1.INIT1 = 16'h5555;
    defparam sub_59_add_2_1.INJECT1_0 = "NO";
    defparam sub_59_add_2_1.INJECT1_1 = "NO";
    LUT4 i14439_2_lut_4_lut (.A(count[8]), .B(n32430), .C(n30563), .D(n925[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14439_2_lut_4_lut.init = 16'h0200;
    LUT4 i14442_2_lut_4_lut (.A(count[8]), .B(n32430), .C(n30563), .D(n925[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14442_2_lut_4_lut.init = 16'h0200;
    LUT4 i14443_2_lut_4_lut (.A(count[8]), .B(n32430), .C(n30563), .D(n925[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14443_2_lut_4_lut.init = 16'h0200;
    LUT4 i14235_2_lut_4_lut (.A(count[8]), .B(n32430), .C(n30563), .D(n925[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i14235_2_lut_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_adj_239 (.A(count[11]), .B(count[10]), .Z(n30465)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_239.init = 16'heeee;
    
endmodule
//
// Verilog Description of module PWMReceiver_U3
//

module PWMReceiver_U3 (debug_c_c, n32341, GND_net, \register[3] , n12138, 
            n31000, n30969, n1009, n28317, rc_ch3_c) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n32341;
    input GND_net;
    output [7:0]\register[3] ;
    input n12138;
    output n31000;
    output n30969;
    output n1009;
    input n28317;
    input rc_ch3_c;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    wire [15:0]n116;
    
    wire n32387, n20320, n32386, n28179, n30497, n152, n103, n154, 
        n14451;
    wire [7:0]n43;
    
    wire n32489, n32496, n32497, n32435, n32498, n30507, n32434, 
        n5, n28468, n28316, n5_adj_126, n30513, n30660, n54, n32385, 
        n10, n1003, n1015, n4, n30404, n4_adj_127, n32452, n16, 
        n26, n30253, n4_adj_128, n32451, n32487, n32413, n30446;
    wire [7:0]n916;
    
    wire n30496, n6, n27341, n27342, n27340, n27339, n27338, n27345, 
        n27344, n27343, n27621, n27620, n27619, n27618;
    
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    LUT4 i24761_3_lut_4_lut_4_lut (.A(n32387), .B(n20320), .C(n32386), 
         .D(n28179), .Z(n30497)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i24761_3_lut_4_lut_4_lut.init = 16'h1110;
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    PFUMX i13410 (.BLUT(n152), .ALUT(n103), .C0(count[3]), .Z(n154));
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_341_4_lut (.A(count[3]), .B(n32489), .C(n32496), 
         .D(n32497), .Z(n32435)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_3_lut_rep_341_4_lut.init = 16'h8000;
    LUT4 i3_3_lut_rep_340_4_lut (.A(count[12]), .B(n32498), .C(n30507), 
         .D(count[13]), .Z(n32434)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_3_lut_rep_340_4_lut.init = 16'hfffe;
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i24732_4_lut (.A(n32498), .B(n5), .C(n28468), .D(n28316), .Z(n31000)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i24732_4_lut.init = 16'h3233;
    LUT4 i1_4_lut (.A(n5_adj_126), .B(n30513), .C(n30660), .D(n20320), 
         .Z(n28316)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccec;
    LUT4 i24701_4_lut (.A(n54), .B(n30513), .C(n32385), .D(n10), .Z(n30969)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i24701_4_lut.init = 16'h3323;
    LUT4 i5_2_lut (.A(n1003), .B(n1015), .Z(n5)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i5_2_lut.init = 16'h4444;
    LUT4 i2_4_lut (.A(count[13]), .B(count[12]), .C(n30507), .D(n4), 
         .Z(n28468)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i1_4_lut_adj_223 (.A(count[9]), .B(count[4]), .C(n30404), .D(n4_adj_127), 
         .Z(n4)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_223.init = 16'hfaea;
    LUT4 i8_4_lut (.A(n32452), .B(n16), .C(count[13]), .D(count[11]), 
         .Z(n14451)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i8_4_lut.init = 16'h0004;
    LUT4 i7_4_lut (.A(count[10]), .B(n32341), .C(n26), .D(n30513), .Z(n16)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i7_4_lut.init = 16'h0040;
    FD1P3IX valid_48 (.D(n30497), .SP(n28317), .CD(GND_net), .CK(debug_c_c), 
            .Q(n1009));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i33_3_lut (.A(n30253), .B(n154), .C(count[9]), .Z(n26)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i33_3_lut.init = 16'h3a3a;
    LUT4 i1_2_lut (.A(n1015), .B(n1003), .Z(n30513)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i2_4_lut_adj_224 (.A(n32496), .B(count[5]), .C(count[3]), .D(n4_adj_128), 
         .Z(n28179)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_4_lut_adj_224.init = 16'h8880;
    LUT4 i1_2_lut_adj_225 (.A(count[11]), .B(count[10]), .Z(n30507)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_225.init = 16'heeee;
    IFS1P3DX latched_in_45 (.D(rc_ch3_c), .SP(n32341), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1015));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_226 (.A(n30404), .B(n32497), .C(count[0]), .D(n32451), 
         .Z(n30253)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_4_lut_adj_226.init = 16'h8000;
    LUT4 i14581_3_lut (.A(count[9]), .B(n32434), .C(n154), .Z(n20320)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i14581_3_lut.init = 16'hecec;
    FD1P3AX prev_in_46 (.D(n1015), .SP(n32341), .CK(debug_c_c), .Q(n1003));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_393 (.A(count[6]), .B(count[7]), .C(count[8]), .Z(n32487)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_393.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut (.A(count[6]), .B(count[7]), .C(count[8]), .D(n32489), 
         .Z(n103)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_319_4_lut (.A(n32452), .B(count[13]), .C(n30507), 
         .D(count[9]), .Z(n32413)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_319_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_227 (.A(n32497), .B(n32496), .C(n32451), .D(count[0]), 
         .Z(n30446)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_227.init = 16'h8000;
    LUT4 i14433_2_lut_4_lut (.A(n32413), .B(count[8]), .C(n32435), .D(n916[7]), 
         .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14433_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_rep_395 (.A(count[4]), .B(count[5]), .Z(n32489)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_rep_395.init = 16'h8888;
    LUT4 i1_2_lut_rep_357_3_lut (.A(count[4]), .B(count[5]), .C(count[3]), 
         .Z(n32451)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_rep_357_3_lut.init = 16'h8080;
    LUT4 i14432_2_lut_4_lut (.A(n32413), .B(count[8]), .C(n32435), .D(n916[6]), 
         .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14432_2_lut_4_lut.init = 16'h0400;
    LUT4 i14431_2_lut_4_lut (.A(n32413), .B(count[8]), .C(n32435), .D(n916[5]), 
         .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14431_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_rep_402 (.A(count[6]), .B(count[7]), .Z(n32496)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_402.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), .Z(n30404)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_403 (.A(count[2]), .B(count[1]), .Z(n32497)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_403.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_228 (.A(count[2]), .B(count[1]), .C(count[4]), 
         .Z(n4_adj_128)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_adj_228.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(count[2]), .B(count[1]), .C(count[5]), .D(count[3]), 
         .Z(n4_adj_127)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_rep_404 (.A(count[15]), .B(count[14]), .Z(n32498)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_404.init = 16'heeee;
    LUT4 i1_2_lut_rep_293_3_lut (.A(count[15]), .B(count[14]), .C(n28468), 
         .Z(n32387)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_293_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_358_3_lut (.A(count[15]), .B(count[14]), .C(count[12]), 
         .Z(n32452)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_358_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[15]), .B(count[14]), .C(n5), .D(n28468), 
         .Z(n30496)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i14430_2_lut_4_lut (.A(n32413), .B(count[8]), .C(n32435), .D(n916[4]), 
         .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14430_2_lut_4_lut.init = 16'h0400;
    LUT4 i14429_2_lut_4_lut (.A(n32413), .B(count[8]), .C(n32435), .D(n916[3]), 
         .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14429_2_lut_4_lut.init = 16'h0400;
    LUT4 i14428_2_lut_4_lut (.A(n32413), .B(count[8]), .C(n32435), .D(n916[2]), 
         .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14428_2_lut_4_lut.init = 16'h0400;
    LUT4 i14427_2_lut_4_lut (.A(n32413), .B(count[8]), .C(n32435), .D(n916[1]), 
         .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14427_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_229 (.A(n32413), .B(count[8]), .C(n32435), 
         .D(n54), .Z(n5_adj_126)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_229.init = 16'h00fb;
    LUT4 i14230_2_lut_4_lut (.A(n32413), .B(count[8]), .C(n32435), .D(n916[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i14230_2_lut_4_lut.init = 16'h0400;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n12138), .PD(n14451), .CK(debug_c_c), 
            .Q(\register[3] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i10_3_lut_3_lut_4_lut (.A(count[8]), .B(n32413), .C(n30446), 
         .D(n28179), .Z(n10)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i10_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_3_lut_rep_291_4_lut (.A(count[9]), .B(n32434), .C(n32435), 
         .D(count[8]), .Z(n32385)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_3_lut_rep_291_4_lut.init = 16'hfeff;
    LUT4 i23_4_lut (.A(n32487), .B(count[2]), .C(n32489), .D(n6), .Z(n152)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'hfaea;
    LUT4 i2_2_lut (.A(count[1]), .B(count[0]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i21_3_lut_4_lut (.A(count[9]), .B(n32434), .C(n20320), .D(n30253), 
         .Z(n54)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i21_3_lut_4_lut.init = 16'h0f0e;
    CCU2D add_1481_9 (.A0(count[7]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27341), 
          .COUT(n27342), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_9.INIT0 = 16'hd222;
    defparam add_1481_9.INIT1 = 16'hd222;
    defparam add_1481_9.INJECT1_0 = "NO";
    defparam add_1481_9.INJECT1_1 = "NO";
    CCU2D add_1481_7 (.A0(count[5]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27340), 
          .COUT(n27341), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_7.INIT0 = 16'hd222;
    defparam add_1481_7.INIT1 = 16'hd222;
    defparam add_1481_7.INJECT1_0 = "NO";
    defparam add_1481_7.INJECT1_1 = "NO";
    CCU2D add_1481_5 (.A0(count[3]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27339), 
          .COUT(n27340), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_5.INIT0 = 16'hd222;
    defparam add_1481_5.INIT1 = 16'hd222;
    defparam add_1481_5.INJECT1_0 = "NO";
    defparam add_1481_5.INJECT1_1 = "NO";
    CCU2D add_1481_3 (.A0(count[1]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27338), 
          .COUT(n27339), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_3.INIT0 = 16'hd222;
    defparam add_1481_3.INIT1 = 16'hd222;
    defparam add_1481_3.INJECT1_0 = "NO";
    defparam add_1481_3.INJECT1_1 = "NO";
    CCU2D add_1481_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n30496), .B1(n1015), .C1(count[0]), .D1(n1003), .COUT(n27338), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_1.INIT0 = 16'hF000;
    defparam add_1481_1.INIT1 = 16'ha565;
    defparam add_1481_1.INJECT1_0 = "NO";
    defparam add_1481_1.INJECT1_1 = "NO";
    LUT4 i24302_3_lut_4_lut (.A(count[8]), .B(n32413), .C(n28179), .D(n30446), 
         .Z(n30660)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i24302_3_lut_4_lut.init = 16'hfeee;
    CCU2D add_1481_17 (.A0(count[15]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27345), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_17.INIT0 = 16'hd222;
    defparam add_1481_17.INIT1 = 16'h0000;
    defparam add_1481_17.INJECT1_0 = "NO";
    defparam add_1481_17.INJECT1_1 = "NO";
    CCU2D add_1481_15 (.A0(count[13]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27344), 
          .COUT(n27345), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_15.INIT0 = 16'hd222;
    defparam add_1481_15.INIT1 = 16'hd222;
    defparam add_1481_15.INJECT1_0 = "NO";
    defparam add_1481_15.INJECT1_1 = "NO";
    CCU2D add_1481_13 (.A0(count[11]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27343), 
          .COUT(n27344), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_13.INIT0 = 16'hd222;
    defparam add_1481_13.INIT1 = 16'hd222;
    defparam add_1481_13.INJECT1_0 = "NO";
    defparam add_1481_13.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27621), 
          .S0(n916[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_58_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_9.INIT1 = 16'h0000;
    defparam sub_58_add_2_9.INJECT1_0 = "NO";
    defparam sub_58_add_2_9.INJECT1_1 = "NO";
    CCU2D add_1481_11 (.A0(count[9]), .B0(n5), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n5), .C1(GND_net), .D1(GND_net), .CIN(n27342), 
          .COUT(n27343), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1481_11.INIT0 = 16'hd222;
    defparam add_1481_11.INIT1 = 16'hd222;
    defparam add_1481_11.INJECT1_0 = "NO";
    defparam add_1481_11.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27620), 
          .COUT(n27621), .S0(n916[5]), .S1(n916[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_58_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_58_add_2_7.INJECT1_0 = "NO";
    defparam sub_58_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27619), 
          .COUT(n27620), .S0(n916[3]), .S1(n916[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_58_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_58_add_2_5.INJECT1_0 = "NO";
    defparam sub_58_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27618), 
          .COUT(n27619), .S0(n916[1]), .S1(n916[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_58_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_58_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_58_add_2_3.INJECT1_0 = "NO";
    defparam sub_58_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_58_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27618), 
          .S1(n916[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_58_add_2_1.INIT0 = 16'hF000;
    defparam sub_58_add_2_1.INIT1 = 16'h5555;
    defparam sub_58_add_2_1.INJECT1_0 = "NO";
    defparam sub_58_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_292_3_lut (.A(count[9]), .B(n32434), .C(count[8]), 
         .Z(n32386)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_292_3_lut.init = 16'hfefe;
    
endmodule
//
// Verilog Description of module PWMReceiver_U4
//

module PWMReceiver_U4 (n1000, n988, n32341, debug_c_c, GND_net, \register[2] , 
            n32336, n14446, n994, rc_ch2_c, n54, n4) /* synthesis syn_module_defined=1 */ ;
    output n1000;
    output n988;
    input n32341;
    input debug_c_c;
    input GND_net;
    output [7:0]\register[2] ;
    input n32336;
    input n14446;
    output n994;
    input rc_ch2_c;
    output n54;
    output n4;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    
    wire n32491, n28253, n4_c, n30443, n28193, n28059, n32471, 
        n4_adj_123, n5, n30654, n20380, n8, n30444, n32333, n30453, 
        n32490;
    wire [15:0]n116;
    wire [7:0]n43;
    
    wire n30367, n29666, n11825, n32519, n63, n21771, n30744, 
        n30520, n32427, n4_adj_124, n30267, n32426, n32447, n25, 
        n11, n6, n27353, n27352, n27351, n27350, n27349, n27348, 
        n27347, n27346, n27625;
    wire [7:0]n907;
    
    wire n27624, n27623, n27622, n29792, n28382, n32520;
    
    LUT4 i1_3_lut_4_lut (.A(count[8]), .B(n32491), .C(count[9]), .D(n28253), 
         .Z(n4_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i24753_4_lut (.A(n1000), .B(n30443), .C(n988), .D(n32341), 
         .Z(n28193)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(D)))) */ ;
    defparam i24753_4_lut.init = 16'h3100;
    LUT4 i1_4_lut (.A(n28059), .B(n32471), .C(n988), .D(n4_adj_123), 
         .Z(n30443)) /* synthesis lut_function=(!(A+(B+!((D)+!C)))) */ ;
    defparam i1_4_lut.init = 16'h1101;
    LUT4 i1_4_lut_adj_204 (.A(n1000), .B(n5), .C(n30654), .D(n20380), 
         .Z(n4_adj_123)) /* synthesis lut_function=(A+!(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_204.init = 16'haaea;
    LUT4 i2_4_lut (.A(n32471), .B(count[12]), .C(n8), .D(count[11]), 
         .Z(n30444)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_4_lut.init = 16'h0010;
    LUT4 i3_3_lut (.A(n32333), .B(count[10]), .C(count[13]), .Z(n8)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i3_3_lut.init = 16'h0202;
    LUT4 i2_4_lut_adj_205 (.A(count[12]), .B(n30453), .C(count[13]), .D(n4_c), 
         .Z(n28059)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_205.init = 16'ha080;
    LUT4 i2_4_lut_adj_206 (.A(count[3]), .B(count[5]), .C(n32490), .D(count[4]), 
         .Z(n28253)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_4_lut_adj_206.init = 16'hffec;
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n32336), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i1_4_lut_else_4_lut (.A(n30367), .B(n29666), .C(n11825), .D(count[9]), 
         .Z(n32519)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h0002;
    FD1P3AX valid_48 (.D(n30444), .SP(n28193), .CK(debug_c_c), .Q(n994));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(n1000), .B(n988), .Z(n63)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_adj_207 (.A(n1000), .B(n988), .Z(n21771)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_adj_207.init = 16'h2222;
    LUT4 count_8__bdd_4_lut (.A(count[8]), .B(n30367), .C(n30744), .D(count[9]), 
         .Z(n32333)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam count_8__bdd_4_lut.init = 16'hf0ee;
    LUT4 i24216_2_lut_rep_377 (.A(count[14]), .B(count[15]), .Z(n32471)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24216_2_lut_rep_377.init = 16'heeee;
    LUT4 i2_3_lut_4_lut (.A(count[14]), .B(count[15]), .C(n21771), .D(n28059), 
         .Z(n30520)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_333 (.A(count[9]), .B(n11825), .Z(n32427)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i1_2_lut_rep_333.init = 16'heeee;
    IFS1P3DX latched_in_45 (.D(rc_ch2_c), .SP(n32341), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n1000));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_396 (.A(count[2]), .B(count[1]), .Z(n32490)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_396.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count[2]), .B(count[1]), .C(count[3]), .Z(n4_adj_124)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_397 (.A(count[6]), .B(count[7]), .Z(n32491)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_397.init = 16'h8888;
    LUT4 i1_2_lut_rep_332_3_lut (.A(count[6]), .B(count[7]), .C(n30267), 
         .Z(n32426)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_332_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count[6]), .B(count[7]), .C(count[0]), 
         .D(n30267), .Z(n29666)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_353_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n32447)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_353_3_lut.init = 16'h8080;
    FD1P3AX prev_in_46 (.D(n1000), .SP(n32341), .CK(debug_c_c), .Q(n988));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n32336), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n32336), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n32336), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n32336), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n32336), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n32336), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n32336), .PD(n14446), .CK(debug_c_c), 
            .Q(\register[2] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    LUT4 i24809_4_lut (.A(count[8]), .B(count[7]), .C(n25), .D(count[6]), 
         .Z(n30744)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i24809_4_lut.init = 16'h0001;
    LUT4 i1_4_lut_adj_208 (.A(count[0]), .B(n11), .C(n6), .D(count[1]), 
         .Z(n25)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_208.init = 16'hccc8;
    LUT4 i2_2_lut (.A(count[3]), .B(count[2]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_209 (.A(n32491), .B(count[5]), .C(count[4]), .D(n4_adj_124), 
         .Z(n30367)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_209.init = 16'h8880;
    LUT4 i1_2_lut_adj_210 (.A(count[5]), .B(count[4]), .Z(n11)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_adj_210.init = 16'h8888;
    CCU2D add_1477_17 (.A0(count[15]), .B0(n63), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27353), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_17.INIT0 = 16'h7888;
    defparam add_1477_17.INIT1 = 16'h0000;
    defparam add_1477_17.INJECT1_0 = "NO";
    defparam add_1477_17.INJECT1_1 = "NO";
    CCU2D add_1477_15 (.A0(n63), .B0(count[13]), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n63), .C1(GND_net), .D1(GND_net), .CIN(n27352), 
          .COUT(n27353), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_15.INIT0 = 16'h7888;
    defparam add_1477_15.INIT1 = 16'h7888;
    defparam add_1477_15.INJECT1_0 = "NO";
    defparam add_1477_15.INJECT1_1 = "NO";
    CCU2D add_1477_13 (.A0(count[11]), .B0(n21771), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n63), .C1(GND_net), .D1(GND_net), .CIN(n27351), 
          .COUT(n27352), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_13.INIT0 = 16'hd222;
    defparam add_1477_13.INIT1 = 16'h7888;
    defparam add_1477_13.INJECT1_0 = "NO";
    defparam add_1477_13.INJECT1_1 = "NO";
    CCU2D add_1477_11 (.A0(count[9]), .B0(n21771), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n21771), .C1(GND_net), .D1(GND_net), .CIN(n27350), 
          .COUT(n27351), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_11.INIT0 = 16'hd222;
    defparam add_1477_11.INIT1 = 16'hd222;
    defparam add_1477_11.INJECT1_0 = "NO";
    defparam add_1477_11.INJECT1_1 = "NO";
    CCU2D add_1477_9 (.A0(count[7]), .B0(n21771), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n21771), .C1(GND_net), .D1(GND_net), .CIN(n27349), 
          .COUT(n27350), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_9.INIT0 = 16'hd222;
    defparam add_1477_9.INIT1 = 16'hd222;
    defparam add_1477_9.INJECT1_0 = "NO";
    defparam add_1477_9.INJECT1_1 = "NO";
    CCU2D add_1477_7 (.A0(count[5]), .B0(n21771), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n21771), .C1(GND_net), .D1(GND_net), .CIN(n27348), 
          .COUT(n27349), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_7.INIT0 = 16'hd222;
    defparam add_1477_7.INIT1 = 16'hd222;
    defparam add_1477_7.INJECT1_0 = "NO";
    defparam add_1477_7.INJECT1_1 = "NO";
    CCU2D add_1477_5 (.A0(count[3]), .B0(n21771), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n21771), .C1(GND_net), .D1(GND_net), .CIN(n27347), 
          .COUT(n27348), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_5.INIT0 = 16'hd222;
    defparam add_1477_5.INIT1 = 16'hd222;
    defparam add_1477_5.INJECT1_0 = "NO";
    defparam add_1477_5.INJECT1_1 = "NO";
    CCU2D add_1477_3 (.A0(count[1]), .B0(n21771), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n21771), .C1(GND_net), .D1(GND_net), .CIN(n27346), 
          .COUT(n27347), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_3.INIT0 = 16'hd222;
    defparam add_1477_3.INIT1 = 16'hd222;
    defparam add_1477_3.INJECT1_0 = "NO";
    defparam add_1477_3.INJECT1_1 = "NO";
    CCU2D add_1477_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n30520), .B1(n1000), .C1(count[0]), .D1(n988), .COUT(n27346), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1477_1.INIT0 = 16'hF000;
    defparam add_1477_1.INIT1 = 16'ha565;
    defparam add_1477_1.INJECT1_0 = "NO";
    defparam add_1477_1.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27625), 
          .S0(n907[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_57_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_9.INIT1 = 16'h0000;
    defparam sub_57_add_2_9.INJECT1_0 = "NO";
    defparam sub_57_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27624), 
          .COUT(n27625), .S0(n907[5]), .S1(n907[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_57_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_57_add_2_7.INJECT1_0 = "NO";
    defparam sub_57_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27623), 
          .COUT(n27624), .S0(n907[3]), .S1(n907[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_57_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_57_add_2_5.INJECT1_0 = "NO";
    defparam sub_57_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27622), 
          .COUT(n27623), .S0(n907[1]), .S1(n907[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_57_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_57_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_57_add_2_3.INJECT1_0 = "NO";
    defparam sub_57_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_57_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27622), 
          .S1(n907[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_57_add_2_1.INIT0 = 16'hF000;
    defparam sub_57_add_2_1.INIT1 = 16'h5555;
    defparam sub_57_add_2_1.INJECT1_0 = "NO";
    defparam sub_57_add_2_1.INJECT1_1 = "NO";
    LUT4 i24298_3_lut_4_lut (.A(count[8]), .B(n32427), .C(n30367), .D(n29666), 
         .Z(n30654)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[28:39])
    defparam i24298_3_lut_4_lut.init = 16'hfeee;
    LUT4 i1_2_lut_4_lut (.A(n32426), .B(count[8]), .C(n32427), .D(n907[0]), 
         .Z(n43[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_211 (.A(n32426), .B(count[8]), .C(n32427), 
         .D(n54), .Z(n5)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_211.init = 16'h00fb;
    LUT4 i1_2_lut_4_lut_adj_212 (.A(n32426), .B(count[8]), .C(n32427), 
         .D(n907[7]), .Z(n43[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_212.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_213 (.A(n32426), .B(count[8]), .C(n32427), 
         .D(n907[6]), .Z(n43[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_213.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_214 (.A(n32426), .B(count[8]), .C(n32427), 
         .D(n907[5]), .Z(n43[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_214.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_215 (.A(n32426), .B(count[8]), .C(n32427), 
         .D(n907[4]), .Z(n43[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_215.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_216 (.A(n32426), .B(count[8]), .C(n32427), 
         .D(n907[3]), .Z(n43[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_216.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_217 (.A(n32426), .B(count[8]), .C(n32427), 
         .D(n907[2]), .Z(n43[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_217.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_218 (.A(n32426), .B(count[8]), .C(n32427), 
         .D(n907[1]), .Z(n43[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_218.init = 16'h0400;
    LUT4 i3_4_lut (.A(count[3]), .B(n11), .C(count[1]), .D(count[2]), 
         .Z(n30267)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i3_4_lut_adj_219 (.A(count[13]), .B(n30453), .C(count[12]), .D(n32471), 
         .Z(n11825)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_219.init = 16'hfffe;
    LUT4 i1_2_lut_adj_220 (.A(count[10]), .B(count[11]), .Z(n30453)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_220.init = 16'heeee;
    LUT4 i21_4_lut (.A(n29792), .B(n20380), .C(n32427), .D(n32447), 
         .Z(n54)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[13:39])
    defparam i21_4_lut.init = 16'h3230;
    LUT4 i1_2_lut_adj_221 (.A(count[0]), .B(n30267), .Z(n29792)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_adj_221.init = 16'h8888;
    LUT4 i14641_3_lut (.A(n28382), .B(n11825), .C(count[9]), .Z(n20380)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i14641_3_lut.init = 16'hecec;
    LUT4 i3_4_lut_adj_222 (.A(n25), .B(count[6]), .C(count[8]), .D(count[7]), 
         .Z(n28382)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_222.init = 16'hfffe;
    LUT4 i1_4_lut_then_4_lut (.A(n32491), .B(n11825), .C(count[9]), .D(n30267), 
         .Z(n32520)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B+(C)))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0103;
    PFUMX i25261 (.BLUT(n32519), .ALUT(n32520), .C0(count[8]), .Z(n4));
    
endmodule
//
// Verilog Description of module PWMReceiver_U5
//

module PWMReceiver_U5 (debug_c_c, n32341, GND_net, \register[1] , n12841, 
            n31049, n979, n28312, rc_ch1_c, n30911) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n32341;
    input GND_net;
    output [7:0]\register[1] ;
    input n12841;
    output n31049;
    output n979;
    input n28312;
    input rc_ch1_c;
    output n30911;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire [15:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    wire [15:0]n116;
    
    wire n14448;
    wire [7:0]n43;
    
    wire n30245, n4, n973, n985, n32474, n32404, n30503, n32477, 
        n28217, n11792, n32428, n32406, n20451, n32405, n30247, 
        n32377, n32378, n30579, n23, n30716, n30502, n27361, n27360, 
        n27359, n27358, n32355, n27357, n27356, n27355, n27354, 
        n27629;
    wire [7:0]n898;
    
    wire n27628, n27627, n27626, n30156, n30437, n30474, n28385, 
        n30476, n6, n95, n11845, n49_adj_122, n30750, n30722;
    
    FD1P3IX count_i0_i0 (.D(n116[0]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i0.GSR = "ENABLED";
    FD1P3JX period_i0_i0 (.D(n43[0]), .SP(n12841), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut (.A(count[6]), .B(count[7]), .C(count[5]), .Z(n30245)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_194 (.A(count[6]), .B(count[7]), .C(count[8]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i1_2_lut_3_lut_adj_194.init = 16'h8080;
    LUT4 i5_2_lut_rep_380 (.A(n973), .B(n985), .Z(n32474)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i5_2_lut_rep_380.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_195 (.A(n973), .B(n985), .C(n32404), .Z(n30503)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(154[10:31])
    defparam i1_2_lut_3_lut_adj_195.init = 16'hf4f4;
    LUT4 i1_2_lut_rep_383 (.A(n985), .B(n973), .Z(n32477)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_383.init = 16'hbbbb;
    LUT4 i24781_2_lut_3_lut (.A(n985), .B(n973), .C(n28217), .Z(n31049)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i24781_2_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_334 (.A(count[9]), .B(n11792), .Z(n32428)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i1_2_lut_rep_334.init = 16'heeee;
    LUT4 i14712_2_lut_3_lut_4_lut (.A(count[9]), .B(n11792), .C(n32406), 
         .D(count[8]), .Z(n20451)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i14712_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_311_3_lut (.A(count[9]), .B(n11792), .C(count[8]), 
         .Z(n32405)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i1_2_lut_rep_311_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_283_3_lut_4_lut (.A(count[9]), .B(n11792), .C(n30247), 
         .D(count[8]), .Z(n32377)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[28:39])
    defparam i1_2_lut_rep_283_3_lut_4_lut.init = 16'hfffe;
    LUT4 i24357_3_lut_4_lut (.A(n32378), .B(n30579), .C(n32428), .D(n23), 
         .Z(n30716)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(172[13:39])
    defparam i24357_3_lut_4_lut.init = 16'hfffe;
    FD1P3AX valid_48 (.D(n30502), .SP(n28312), .CK(debug_c_c), .Q(n979));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam valid_48.GSR = "ENABLED";
    FD1P3IX count_i0_i15 (.D(n116[15]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i15.GSR = "ENABLED";
    FD1P3IX count_i0_i14 (.D(n116[14]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i14.GSR = "ENABLED";
    FD1P3JX count_i0_i13 (.D(n116[13]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i13.GSR = "ENABLED";
    FD1P3JX count_i0_i12 (.D(n116[12]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i12.GSR = "ENABLED";
    FD1P3IX count_i0_i11 (.D(n116[11]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i11.GSR = "ENABLED";
    FD1P3IX count_i0_i10 (.D(n116[10]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i10.GSR = "ENABLED";
    FD1P3IX count_i0_i9 (.D(n116[9]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i9.GSR = "ENABLED";
    FD1P3JX count_i0_i8 (.D(n116[8]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i8.GSR = "ENABLED";
    FD1P3JX count_i0_i7 (.D(n116[7]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i7.GSR = "ENABLED";
    FD1P3AX prev_in_46 (.D(n985), .SP(n32341), .CK(debug_c_c), .Q(n973));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam prev_in_46.GSR = "ENABLED";
    FD1P3JX count_i0_i6 (.D(n116[6]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i6.GSR = "ENABLED";
    IFS1P3DX latched_in_45 (.D(rc_ch1_c), .SP(n32341), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(n985));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam latched_in_45.GSR = "ENABLED";
    FD1P3IX count_i0_i5 (.D(n116[5]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i5.GSR = "ENABLED";
    FD1P3IX count_i0_i4 (.D(n116[4]), .SP(n32341), .CD(GND_net), .CK(debug_c_c), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i4.GSR = "ENABLED";
    FD1P3JX count_i0_i3 (.D(n116[3]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i3.GSR = "ENABLED";
    FD1P3JX count_i0_i2 (.D(n116[2]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i2.GSR = "ENABLED";
    FD1P3JX count_i0_i1 (.D(n116[1]), .SP(n32341), .PD(GND_net), .CK(debug_c_c), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam count_i0_i1.GSR = "ENABLED";
    FD1P3JX period_i0_i7 (.D(n43[7]), .SP(n12841), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i7.GSR = "ENABLED";
    FD1P3JX period_i0_i6 (.D(n43[6]), .SP(n12841), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i6.GSR = "ENABLED";
    FD1P3JX period_i0_i5 (.D(n43[5]), .SP(n12841), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i5.GSR = "ENABLED";
    FD1P3JX period_i0_i4 (.D(n43[4]), .SP(n12841), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i4.GSR = "ENABLED";
    FD1P3JX period_i0_i3 (.D(n43[3]), .SP(n12841), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i3.GSR = "ENABLED";
    FD1P3JX period_i0_i2 (.D(n43[2]), .SP(n12841), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i2.GSR = "ENABLED";
    FD1P3JX period_i0_i1 (.D(n43[1]), .SP(n12841), .PD(n14448), .CK(debug_c_c), 
            .Q(\register[1] [1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam period_i0_i1.GSR = "ENABLED";
    CCU2D add_1473_17 (.A0(count[15]), .B0(n32474), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27361), 
          .S0(n116[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_17.INIT0 = 16'hd222;
    defparam add_1473_17.INIT1 = 16'h0000;
    defparam add_1473_17.INJECT1_0 = "NO";
    defparam add_1473_17.INJECT1_1 = "NO";
    CCU2D add_1473_15 (.A0(count[13]), .B0(n32474), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(n32474), .C1(GND_net), .D1(GND_net), .CIN(n27360), 
          .COUT(n27361), .S0(n116[13]), .S1(n116[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_15.INIT0 = 16'hd222;
    defparam add_1473_15.INIT1 = 16'hd222;
    defparam add_1473_15.INJECT1_0 = "NO";
    defparam add_1473_15.INJECT1_1 = "NO";
    CCU2D add_1473_13 (.A0(count[11]), .B0(n32474), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(n32474), .C1(GND_net), .D1(GND_net), .CIN(n27359), 
          .COUT(n27360), .S0(n116[11]), .S1(n116[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_13.INIT0 = 16'hd222;
    defparam add_1473_13.INIT1 = 16'hd222;
    defparam add_1473_13.INJECT1_0 = "NO";
    defparam add_1473_13.INJECT1_1 = "NO";
    CCU2D add_1473_11 (.A0(count[9]), .B0(n32474), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(n32474), .C1(GND_net), .D1(GND_net), .CIN(n27358), 
          .COUT(n27359), .S0(n116[9]), .S1(n116[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_11.INIT0 = 16'hd222;
    defparam add_1473_11.INIT1 = 16'hd222;
    defparam add_1473_11.INJECT1_0 = "NO";
    defparam add_1473_11.INJECT1_1 = "NO";
    LUT4 i21_3_lut_rep_261_4_lut (.A(count[8]), .B(n32406), .C(n32428), 
         .D(n30579), .Z(n32355)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i21_3_lut_rep_261_4_lut.init = 16'h00f8;
    CCU2D add_1473_9 (.A0(count[7]), .B0(n32474), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(n32474), .C1(GND_net), .D1(GND_net), .CIN(n27357), 
          .COUT(n27358), .S0(n116[7]), .S1(n116[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_9.INIT0 = 16'hd222;
    defparam add_1473_9.INIT1 = 16'hd222;
    defparam add_1473_9.INJECT1_0 = "NO";
    defparam add_1473_9.INJECT1_1 = "NO";
    CCU2D add_1473_7 (.A0(count[5]), .B0(n32474), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(n32474), .C1(GND_net), .D1(GND_net), .CIN(n27356), 
          .COUT(n27357), .S0(n116[5]), .S1(n116[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_7.INIT0 = 16'hd222;
    defparam add_1473_7.INIT1 = 16'hd222;
    defparam add_1473_7.INJECT1_0 = "NO";
    defparam add_1473_7.INJECT1_1 = "NO";
    CCU2D add_1473_5 (.A0(count[3]), .B0(n32474), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(n32474), .C1(GND_net), .D1(GND_net), .CIN(n27355), 
          .COUT(n27356), .S0(n116[3]), .S1(n116[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_5.INIT0 = 16'hd222;
    defparam add_1473_5.INIT1 = 16'hd222;
    defparam add_1473_5.INJECT1_0 = "NO";
    defparam add_1473_5.INJECT1_1 = "NO";
    CCU2D add_1473_3 (.A0(count[1]), .B0(n32474), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(n32474), .C1(GND_net), .D1(GND_net), .CIN(n27354), 
          .COUT(n27355), .S0(n116[1]), .S1(n116[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_3.INIT0 = 16'hd222;
    defparam add_1473_3.INIT1 = 16'hd222;
    defparam add_1473_3.INJECT1_0 = "NO";
    defparam add_1473_3.INJECT1_1 = "NO";
    CCU2D add_1473_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n30503), .B1(n985), .C1(count[0]), .D1(n973), .COUT(n27354), 
          .S1(n116[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(159[7] 186[10])
    defparam add_1473_1.INIT0 = 16'hF000;
    defparam add_1473_1.INIT1 = 16'ha565;
    defparam add_1473_1.INJECT1_0 = "NO";
    defparam add_1473_1.INJECT1_1 = "NO";
    CCU2D sub_56_add_2_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27629), 
          .S0(n898[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_56_add_2_9.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_9.INIT1 = 16'h0000;
    defparam sub_56_add_2_9.INJECT1_0 = "NO";
    defparam sub_56_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_56_add_2_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27628), 
          .COUT(n27629), .S0(n898[5]), .S1(n898[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_56_add_2_7.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_7.INIT1 = 16'h5aaa;
    defparam sub_56_add_2_7.INJECT1_0 = "NO";
    defparam sub_56_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_56_add_2_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27627), 
          .COUT(n27628), .S0(n898[3]), .S1(n898[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_56_add_2_5.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_5.INIT1 = 16'h5aaa;
    defparam sub_56_add_2_5.INJECT1_0 = "NO";
    defparam sub_56_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_56_add_2_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27626), 
          .COUT(n27627), .S0(n898[1]), .S1(n898[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_56_add_2_3.INIT0 = 16'h5aaa;
    defparam sub_56_add_2_3.INIT1 = 16'h5aaa;
    defparam sub_56_add_2_3.INJECT1_0 = "NO";
    defparam sub_56_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_56_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27626), 
          .S1(n898[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(170[22:33])
    defparam sub_56_add_2_1.INIT0 = 16'hF000;
    defparam sub_56_add_2_1.INIT1 = 16'h5555;
    defparam sub_56_add_2_1.INJECT1_0 = "NO";
    defparam sub_56_add_2_1.INJECT1_1 = "NO";
    LUT4 i3_4_lut (.A(n973), .B(n32341), .C(n30156), .D(n30579), .Z(n14448)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut.init = 16'h0080;
    LUT4 i2_4_lut (.A(n32378), .B(n28217), .C(count[9]), .D(n985), .Z(n30156)) /* synthesis lut_function=(!(A ((D)+!B)+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i2_4_lut.init = 16'h00c8;
    LUT4 i14222_2_lut (.A(n898[0]), .B(n23), .Z(n43[0])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14222_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_196 (.A(n32355), .B(n23), .C(n32377), .D(n20451), 
         .Z(n28217)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i2_4_lut_adj_196.init = 16'heefe;
    LUT4 i24643_4_lut (.A(n30437), .B(n32474), .C(n32404), .D(n32477), 
         .Z(n30911)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i24643_4_lut.init = 16'h3031;
    LUT4 i3_4_lut_adj_197 (.A(n32405), .B(n30716), .C(n32406), .D(n30247), 
         .Z(n30437)) /* synthesis lut_function=(!(A (B)+!A (B+!(C (D))))) */ ;
    defparam i3_4_lut_adj_197.init = 16'h3222;
    LUT4 i2_4_lut_adj_198 (.A(n30474), .B(count[9]), .C(n28385), .D(n4), 
         .Z(n30476)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_198.init = 16'hfeee;
    LUT4 i2_4_lut_adj_199 (.A(count[5]), .B(count[4]), .C(n6), .D(count[3]), 
         .Z(n28385)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(135[16:21])
    defparam i2_4_lut_adj_199.init = 16'hfeee;
    LUT4 i3_4_lut_adj_200 (.A(count[3]), .B(count[4]), .C(count[2]), .D(n30245), 
         .Z(n95)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i3_4_lut_adj_200.init = 16'h8000;
    LUT4 i3_4_lut_adj_201 (.A(count[12]), .B(count[13]), .C(n11845), .D(n30474), 
         .Z(n11792)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_201.init = 16'hfffe;
    LUT4 i1_2_lut (.A(count[15]), .B(count[14]), .Z(n11845)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_202 (.A(count[11]), .B(count[10]), .Z(n30474)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_202.init = 16'heeee;
    LUT4 i1_4_lut (.A(count[8]), .B(n32428), .C(count[1]), .D(n95), 
         .Z(n23)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0222;
    LUT4 i24224_4_lut (.A(n11792), .B(count[9]), .C(n49_adj_122), .D(n30750), 
         .Z(n30579)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i24224_4_lut.init = 16'heeea;
    LUT4 i2_3_lut (.A(count[6]), .B(count[7]), .C(count[8]), .Z(n49_adj_122)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i24391_4_lut (.A(count[4]), .B(count[1]), .C(count[5]), .D(n30722), 
         .Z(n30750)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i24391_4_lut.init = 16'ha080;
    LUT4 i24363_3_lut (.A(count[0]), .B(count[2]), .C(count[3]), .Z(n30722)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i24363_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_203 (.A(count[4]), .B(n30245), .C(count[3]), .D(n6), 
         .Z(n30247)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_4_lut_adj_203.init = 16'hccc8;
    LUT4 i2786_2_lut (.A(count[1]), .B(count[2]), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2786_2_lut.init = 16'h8888;
    LUT4 i24650_3_lut_4_lut_4_lut (.A(n32404), .B(n30579), .C(n32405), 
         .D(n30247), .Z(n30502)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i24650_3_lut_4_lut_4_lut.init = 16'h1110;
    LUT4 i24207_4_lut_rep_310 (.A(n11845), .B(count[13]), .C(count[12]), 
         .D(n30476), .Z(n32404)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i24207_4_lut_rep_310.init = 16'heaaa;
    LUT4 i2_3_lut_rep_312 (.A(n95), .B(count[1]), .C(count[0]), .Z(n32406)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i2_3_lut_rep_312.init = 16'h8080;
    LUT4 i1_2_lut_rep_284_4_lut (.A(n95), .B(count[1]), .C(count[0]), 
         .D(count[8]), .Z(n32378)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(139[9] 188[6])
    defparam i1_2_lut_rep_284_4_lut.init = 16'h8000;
    LUT4 i14426_2_lut (.A(n898[7]), .B(n23), .Z(n43[7])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14426_2_lut.init = 16'h8888;
    LUT4 i14425_2_lut (.A(n898[6]), .B(n23), .Z(n43[6])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14425_2_lut.init = 16'h8888;
    LUT4 i14424_2_lut (.A(n898[5]), .B(n23), .Z(n43[5])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14424_2_lut.init = 16'h8888;
    LUT4 i14423_2_lut (.A(n898[4]), .B(n23), .Z(n43[4])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14423_2_lut.init = 16'h8888;
    LUT4 i14422_2_lut (.A(n898[3]), .B(n23), .Z(n43[3])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14422_2_lut.init = 16'h8888;
    LUT4 i14421_2_lut (.A(n898[2]), .B(n23), .Z(n43[2])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14421_2_lut.init = 16'h8888;
    LUT4 i14420_2_lut (.A(n898[1]), .B(n23), .Z(n43[1])) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/pwm.v(167[10] 171[14])
    defparam i14420_2_lut.init = 16'h8888;
    
endmodule
//
// Verilog Description of module \ProtocolInterface(baud_div=12) 
//

module \ProtocolInterface(baud_div=12)  (debug_c_c, register_addr, n32389, 
            n30258, n3363, n30423, n32348, n1318, n1304, n1310, 
            n12098, databus_out, n32444, n32358, databus, n224, 
            n3181, \select[1] , n12788, \sendcount[1] , debug_c_7, 
            \select[2] , \select[4] , \select[7] , \steps_reg[4] , n15, 
            n9, n30310, n32343, n224_adj_42, n3451, \steps_reg[7] , 
            n13, \steps_reg[3] , n15_adj_33, rw, \steps_reg[5] , n14, 
            n4, n34317, \steps_reg[5]_adj_34 , n14_adj_35, \steps_reg[3]_adj_36 , 
            n15_adj_37, \steps_reg[5]_adj_38 , n14_adj_39, \steps_reg[3]_adj_40 , 
            n15_adj_41, n32513, n11271, n5, n6, \reg_size[2] , n32486, 
            debug_c_2, debug_c_3, debug_c_4, debug_c_5, n34320, n32503, 
            n30401, n11753, \reset_count[14] , \reset_count[12] , \reset_count[13] , 
            \reset_count[11] , n19877, \reset_count[8] , n27962, n9395, 
            \reset_count[10] , \reset_count[9] , GND_net, state, n32, 
            \rdata[0] , bclk, n29158, \rdata[1] , n9396_c, n31442, 
            n183, n31427, n32432, n32409, n32495, n32494) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    output [7:0]register_addr;
    input n32389;
    input n30258;
    output n3363;
    input n30423;
    output n32348;
    output n1318;
    output n1304;
    output n1310;
    input n12098;
    output [31:0]databus_out;
    output n32444;
    input n32358;
    input [31:0]databus;
    input [31:0]n224;
    output [31:0]n3181;
    output \select[1] ;
    input n12788;
    output \sendcount[1] ;
    output debug_c_7;
    output \select[2] ;
    output \select[4] ;
    output \select[7] ;
    input \steps_reg[4] ;
    output n15;
    output n9;
    input n30310;
    input n32343;
    input [31:0]n224_adj_42;
    output [31:0]n3451;
    input \steps_reg[7] ;
    output n13;
    input \steps_reg[3] ;
    output n15_adj_33;
    output rw;
    input \steps_reg[5] ;
    output n14;
    output n4;
    output n34317;
    input \steps_reg[5]_adj_34 ;
    output n14_adj_35;
    input \steps_reg[3]_adj_36 ;
    output n15_adj_37;
    input \steps_reg[5]_adj_38 ;
    output n14_adj_39;
    input \steps_reg[3]_adj_40 ;
    output n15_adj_41;
    output n32513;
    input n11271;
    input n5;
    input n6;
    input \reg_size[2] ;
    input n32486;
    output debug_c_2;
    output debug_c_3;
    output debug_c_4;
    output debug_c_5;
    input n34320;
    input n32503;
    input n30401;
    output n11753;
    input \reset_count[14] ;
    input \reset_count[12] ;
    input \reset_count[13] ;
    input \reset_count[11] ;
    output n19877;
    input \reset_count[8] ;
    input n27962;
    output n9395;
    input \reset_count[10] ;
    input \reset_count[9] ;
    input GND_net;
    output [5:0]state;
    output n32;
    output \rdata[0] ;
    output bclk;
    input n29158;
    output \rdata[1] ;
    input n9396_c;
    input n31442;
    input n183;
    input n31427;
    input n32432;
    input n32409;
    input n32495;
    input n32494;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire \select[7]  /* synthesis SET_AS_NETWORK=select[7] */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(462[15:21])
    wire [3:0]bufcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(46[12:20])
    
    wire n32395, n32548, n34314, n14083;
    wire [7:0]tx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(52[12:19])
    
    wire n32421;
    wire [7:0]n2028;
    
    wire n2539;
    wire [7:0]\buffer[1] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n32468;
    wire [7:0]\buffer[0] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]rx_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(50[13:20])
    
    wire n11, n11_adj_10, n11_adj_11, n11_adj_12, n11_adj_13, n11_adj_14, 
        n11_adj_15, n11_adj_16, n11_adj_17, n11_adj_18, n11_adj_19;
    wire [4:0]sendcount;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(54[12:21])
    
    wire n32407, n32380, n20282, n11_adj_20, n11_adj_21, n11_adj_22, 
        n11936;
    wire [7:0]\buffer[2] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n12022, n28243, n34319, n28238, n28252, n28235, n28255, 
        n29192, n29190, n29174, n29154, n29264, n29150, n29196, 
        n29200, n29152, n29260, n29262, n29266, n29326, n29198, 
        n29186, n11_adj_23, n11_adj_24, n30278, n29727;
    wire [31:0]n1286;
    
    wire n10677, n9437, n29350, n10675, n9441, n1398, n1397, n1391, 
        n30166, n30109, n10751, n29412, n29464, n29726, n13424;
    wire [7:0]esc_data;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(51[12:20])
    
    wire n32272, n2541, n32515, n32461, n4_c, n32545;
    wire [7:0]n9241;
    
    wire n4_adj_25, n32542, n4_adj_26, n32533, n29188, busy, n14425, 
        n29730, n32523;
    wire [7:0]\buffer[3] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n32522, n35, n30114, n6_c, n11639, n1687, escape, n13_c, 
        n11539, n32526, n32525, n32529, n29974, n32528, n30619, 
        n31474, n30106, n15_c, n30714, n32532, n11477, n29621, 
        n14082, n32531, n2497, n30279, n14122, n9_c, n32464;
    wire [4:0]n18;
    
    wire n32535, n32534;
    wire [4:0]n19;
    
    wire n31398, n32476, n32536, n32270, n32271, n4_adj_28, n32524, 
        n32463, n8, n13423, n32538, n4_adj_29, n32527, n4_adj_30, 
        n32530, n4_adj_31, n32539, n32537, n32541, n32540, n32469, 
        n32445, n28389, n32544, n8679, n32543, n32547, n32546, 
        n33741, n33743;
    wire [3:0]n8204;
    wire [7:0]\buffer[4] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    wire [7:0]\buffer[5] ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(45[12:18])
    
    wire n32462;
    wire [3:0]n1682;
    
    wire n9337, n30754, n30175, n30179, n30184, n30177, n30183, 
        n14_adj_43, n30182, n30487, n30185, n30488, n30186, n7, 
        n32470, n30187, n30188, n30189, n30193, n30512, n30178, 
        n30511, n30192, n30194, n30191, n30190, n30181, n30195, 
        n30196, n5_c, n28336, n30198, n30180, n30197, n30201, 
        n32475, n30200, n30176, n28153, n30202, n17, n31399, n30203, 
        n30204, n30206, n30199, n30205, n32478, n5_adj_50, n28343, 
        n30537, n55, n32266, n32482, n32483, n9_adj_53, n32484, 
        n8_adj_57, n5_adj_58, n28341, n18427, n6_adj_59, send, n28369, 
        n11238, n32516, n32517, n5_adj_61, n10, n30705, n30, n31947, 
        n31948, n5_adj_65, n28338, n5_adj_69, n28305, n5_adj_70, 
        n28358, n5_adj_71, n28370;
    wire [7:0]n4846;
    
    wire n7986, n28240, n28251, n28228, n28323, n28306, n28197, 
        n28223, n28297, n28200, n28206, n28201, n28204, n28190, 
        n28344, n28184, n28314, n28283, n28339, n28303, n28302, 
        n5_adj_72, n6_adj_73, n5_adj_74, n5_adj_75, n5_adj_80, n5_adj_81, 
        n5_adj_86, n5_adj_88, n1, n6_adj_91, n8_adj_95, n4_adj_96, 
        n6_adj_97, n6_adj_98, n30390, n5_adj_100, n5_adj_101, n5_adj_102, 
        n5_adj_103, n5_adj_104, n5_adj_105, n5_adj_106, n30734, n5_adj_108, 
        n30708, n5_adj_109, n5_adj_110, n5_adj_111, n5_adj_112, n5_adj_114, 
        n5_adj_115, n5_adj_116, n38, n8_adj_117, n5_adj_118, n5_adj_119;
    
    FD1S3IX bufcount__i3 (.D(n32548), .CK(debug_c_c), .CD(n32395), .Q(bufcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i3.GSR = "ENABLED";
    FD1S3IX bufcount__i2 (.D(n34314), .CK(debug_c_c), .CD(n32395), .Q(bufcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i2.GSR = "ENABLED";
    FD1S3IX bufcount__i1 (.D(n14083), .CK(debug_c_c), .CD(n32395), .Q(bufcount[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i1.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i4 (.D(n2028[4]), .SP(n32421), .CK(debug_c_c), 
            .Q(tx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i3 (.D(n2028[3]), .SP(n32421), .CK(debug_c_c), 
            .Q(tx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i1 (.D(n2028[1]), .SP(n32421), .CK(debug_c_c), 
            .Q(tx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i1.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i7 (.D(\buffer[1] [7]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i7.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut (.A(register_addr[5]), .B(n32389), .C(n30258), 
         .D(register_addr[4]), .Z(n3363)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_3_lut_4_lut.init = 16'h4000;
    LUT4 i2_3_lut_rep_254_4_lut (.A(register_addr[5]), .B(n32389), .C(register_addr[4]), 
         .D(n30423), .Z(n32348)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_3_lut_rep_254_4_lut.init = 16'h4000;
    LUT4 i24_3_lut_4_lut (.A(bufcount[0]), .B(n32468), .C(\buffer[0] [7]), 
         .D(rx_data[7]), .Z(n11)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_52 (.A(bufcount[0]), .B(n32468), .C(\buffer[0] [6]), 
         .D(rx_data[6]), .Z(n11_adj_10)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_52.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_53 (.A(bufcount[0]), .B(n32468), .C(rx_data[5]), 
         .D(\buffer[0] [5]), .Z(n11_adj_11)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_53.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_54 (.A(bufcount[0]), .B(n32468), .C(rx_data[4]), 
         .D(\buffer[0] [4]), .Z(n11_adj_12)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_54.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_55 (.A(bufcount[0]), .B(n32468), .C(rx_data[3]), 
         .D(\buffer[0] [3]), .Z(n11_adj_13)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_55.init = 16'hfe10;
    LUT4 i24_3_lut_4_lut_adj_56 (.A(bufcount[0]), .B(n32468), .C(\buffer[0] [2]), 
         .D(rx_data[2]), .Z(n11_adj_14)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_56.init = 16'hf1e0;
    FD1P3AX reg_addr_i0_i6 (.D(\buffer[1] [6]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i6.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i5 (.D(\buffer[1] [5]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i5.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i4 (.D(\buffer[1] [4]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i4.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i3 (.D(\buffer[1] [3]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i3.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i2 (.D(\buffer[1] [2]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i2.GSR = "ENABLED";
    FD1P3AX reg_addr_i0_i1 (.D(\buffer[1] [1]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i1.GSR = "ENABLED";
    LUT4 i24_3_lut_4_lut_adj_57 (.A(bufcount[0]), .B(n32468), .C(\buffer[0] [1]), 
         .D(rx_data[1]), .Z(n11_adj_15)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_57.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_58 (.A(bufcount[0]), .B(n32468), .C(\buffer[0] [0]), 
         .D(rx_data[0]), .Z(n11_adj_16)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_58.init = 16'hf1e0;
    LUT4 i24_3_lut_4_lut_adj_59 (.A(bufcount[0]), .B(n32468), .C(\buffer[1] [7]), 
         .D(rx_data[7]), .Z(n11_adj_17)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_59.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_60 (.A(bufcount[0]), .B(n32468), .C(\buffer[1] [6]), 
         .D(rx_data[6]), .Z(n11_adj_18)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_60.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_61 (.A(bufcount[0]), .B(n32468), .C(\buffer[1] [5]), 
         .D(rx_data[5]), .Z(n11_adj_19)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_61.init = 16'hf2d0;
    FD1P3IX sendcount__i0 (.D(n20282), .SP(n32407), .CD(n32380), .CK(debug_c_c), 
            .Q(sendcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i0.GSR = "ENABLED";
    LUT4 i24_3_lut_4_lut_adj_62 (.A(bufcount[0]), .B(n32468), .C(\buffer[1] [4]), 
         .D(rx_data[4]), .Z(n11_adj_20)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_62.init = 16'hf2d0;
    LUT4 i24_3_lut_4_lut_adj_63 (.A(bufcount[0]), .B(n32468), .C(rx_data[3]), 
         .D(\buffer[1] [3]), .Z(n11_adj_21)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_63.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_64 (.A(bufcount[0]), .B(n32468), .C(\buffer[1] [2]), 
         .D(rx_data[2]), .Z(n11_adj_22)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_64.init = 16'hf2d0;
    FD1S3JX state_FSM_i1 (.D(n11936), .CK(debug_c_c), .PD(n32395), .Q(n1318));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i1.GSR = "ENABLED";
    FD1P3IX buffer_0___i21 (.D(n28243), .SP(n12022), .CD(n32395), .CK(debug_c_c), 
            .Q(\buffer[2] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i21.GSR = "ENABLED";
    FD1P3IX buffer_0___i20 (.D(n28238), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[2] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i20.GSR = "ENABLED";
    FD1P3IX buffer_0___i19 (.D(n28252), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i19.GSR = "ENABLED";
    FD1P3IX buffer_0___i18 (.D(n28235), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i18.GSR = "ENABLED";
    FD1P3IX buffer_0___i17 (.D(n28255), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i17.GSR = "ENABLED";
    FD1P3IX buffer_0___i16 (.D(n29192), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[1] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i16.GSR = "ENABLED";
    FD1P3IX buffer_0___i15 (.D(n29190), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[1] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i15.GSR = "ENABLED";
    FD1P3IX buffer_0___i14 (.D(n29174), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[1] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i14.GSR = "ENABLED";
    FD1P3IX buffer_0___i13 (.D(n29154), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[1] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i13.GSR = "ENABLED";
    FD1P3IX buffer_0___i12 (.D(n29264), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[1] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i12.GSR = "ENABLED";
    FD1P3IX buffer_0___i11 (.D(n29150), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[1] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i11.GSR = "ENABLED";
    FD1P3IX buffer_0___i10 (.D(n29196), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[1] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i10.GSR = "ENABLED";
    FD1P3IX buffer_0___i9 (.D(n29200), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[1] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i9.GSR = "ENABLED";
    FD1P3IX buffer_0___i8 (.D(n29152), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[0] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i8.GSR = "ENABLED";
    FD1P3IX buffer_0___i7 (.D(n29260), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[0] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i7.GSR = "ENABLED";
    FD1P3IX buffer_0___i6 (.D(n29262), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[0] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i6.GSR = "ENABLED";
    FD1P3IX buffer_0___i5 (.D(n29266), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[0] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i5.GSR = "ENABLED";
    FD1P3IX buffer_0___i4 (.D(n29326), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[0] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i4.GSR = "ENABLED";
    FD1P3IX buffer_0___i3 (.D(n29198), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[0] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i3.GSR = "ENABLED";
    FD1P3IX buffer_0___i2 (.D(n29186), .SP(n12022), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[0] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i2.GSR = "ENABLED";
    LUT4 i24_3_lut_4_lut_adj_65 (.A(bufcount[0]), .B(n32468), .C(rx_data[1]), 
         .D(\buffer[1] [1]), .Z(n11_adj_23)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_65.init = 16'hfd20;
    LUT4 i24_3_lut_4_lut_adj_66 (.A(bufcount[0]), .B(n32468), .C(rx_data[0]), 
         .D(\buffer[1] [0]), .Z(n11_adj_24)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i24_3_lut_4_lut_adj_66.init = 16'hfd20;
    LUT4 i2_3_lut_4_lut (.A(\buffer[0] [0]), .B(n30278), .C(\buffer[0] [2]), 
         .D(\buffer[0] [1]), .Z(n29727)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0400;
    FD1S3IX state_FSM_i21 (.D(n10677), .CK(debug_c_c), .CD(n34319), .Q(n1286[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i21.GSR = "ENABLED";
    FD1S3IX state_FSM_i20 (.D(n9437), .CK(debug_c_c), .CD(n34319), .Q(n1286[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i20.GSR = "ENABLED";
    FD1S3IX state_FSM_i19 (.D(n29350), .CK(debug_c_c), .CD(n32395), .Q(n1286[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i19.GSR = "ENABLED";
    FD1S3IX state_FSM_i18 (.D(n10675), .CK(debug_c_c), .CD(n32395), .Q(n1286[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i18.GSR = "ENABLED";
    FD1S3IX state_FSM_i17 (.D(n9441), .CK(debug_c_c), .CD(n32395), .Q(n1286[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i17.GSR = "ENABLED";
    FD1S3IX state_FSM_i16 (.D(n1398), .CK(debug_c_c), .CD(n32395), .Q(n1286[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i16.GSR = "ENABLED";
    FD1S3IX state_FSM_i15 (.D(n1397), .CK(debug_c_c), .CD(n32395), .Q(n1304));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i15.GSR = "ENABLED";
    FD1S3IX state_FSM_i14 (.D(n1286[12]), .CK(debug_c_c), .CD(n32395), 
            .Q(n1286[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i14.GSR = "ENABLED";
    FD1S3IX state_FSM_i13 (.D(n1286[11]), .CK(debug_c_c), .CD(n32395), 
            .Q(n1286[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i13.GSR = "ENABLED";
    FD1S3IX state_FSM_i12 (.D(n1286[10]), .CK(debug_c_c), .CD(n32395), 
            .Q(n1286[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i12.GSR = "ENABLED";
    FD1S3IX state_FSM_i11 (.D(n1391), .CK(debug_c_c), .CD(n32395), .Q(n1286[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i11.GSR = "ENABLED";
    FD1S3IX state_FSM_i10 (.D(n1310), .CK(debug_c_c), .CD(n32395), .Q(n1286[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i10.GSR = "ENABLED";
    FD1S3IX state_FSM_i9 (.D(n1286[7]), .CK(debug_c_c), .CD(n32395), .Q(n1310));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i9.GSR = "ENABLED";
    FD1S3IX state_FSM_i8 (.D(n1286[6]), .CK(debug_c_c), .CD(n32395), .Q(n1286[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i8.GSR = "ENABLED";
    FD1S3IX state_FSM_i7 (.D(n1286[5]), .CK(debug_c_c), .CD(n32395), .Q(n1286[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i7.GSR = "ENABLED";
    FD1S3IX state_FSM_i6 (.D(n30166), .CK(debug_c_c), .CD(n32395), .Q(n1286[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i6.GSR = "ENABLED";
    FD1S3IX state_FSM_i5 (.D(n30109), .CK(debug_c_c), .CD(n32395), .Q(n1286[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i5.GSR = "ENABLED";
    FD1S3IX state_FSM_i4 (.D(n10751), .CK(debug_c_c), .CD(n32395), .Q(n1286[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i4.GSR = "ENABLED";
    FD1S3IX state_FSM_i3 (.D(n29412), .CK(debug_c_c), .CD(n32395), .Q(n1286[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i3.GSR = "ENABLED";
    FD1S3IX state_FSM_i2 (.D(n29464), .CK(debug_c_c), .CD(n32395), .Q(n1286[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam state_FSM_i2.GSR = "ENABLED";
    LUT4 i2_3_lut_4_lut_adj_67 (.A(\buffer[0] [0]), .B(n30278), .C(\buffer[0] [1]), 
         .D(\buffer[0] [2]), .Z(n29726)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_4_lut_adj_67.init = 16'h0400;
    FD1P3AX reg_addr_i0_i0 (.D(\buffer[1] [0]), .SP(n2539), .CK(debug_c_c), 
            .Q(register_addr[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam reg_addr_i0_i0.GSR = "ENABLED";
    FD1P3AX tx_data_i0_i0 (.D(n2028[0]), .SP(n32421), .CK(debug_c_c), 
            .Q(tx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i0.GSR = "ENABLED";
    FD1S3IX bufcount__i0 (.D(n13424), .CK(debug_c_c), .CD(n32395), .Q(bufcount[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam bufcount__i0.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i0 (.D(n32272), .SP(n12098), .CK(debug_c_c), .Q(esc_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i0.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i0 (.D(\buffer[2] [0]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i0.GSR = "ENABLED";
    LUT4 i882_3_lut (.A(n1286[5]), .B(n32444), .C(n1286[10]), .Z(n2539)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i882_3_lut.init = 16'hc8c8;
    LUT4 mux_429_Mux_1_i7_4_lut_4_lut (.A(n32515), .B(n32461), .C(n4_c), 
         .D(n32545), .Z(n9241[1])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_1_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_2_i7_4_lut_4_lut (.A(n32515), .B(n32461), .C(n4_adj_25), 
         .D(n32542), .Z(n9241[2])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_2_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_4_i7_4_lut_4_lut (.A(n32515), .B(n32461), .C(n4_adj_26), 
         .D(n32533), .Z(n9241[4])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_4_i7_4_lut_4_lut.init = 16'hdc10;
    FD1P3IX buffer_0___i1 (.D(n29188), .SP(n12022), .CD(n32395), .CK(debug_c_c), 
            .Q(\buffer[0] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i1.GSR = "ENABLED";
    LUT4 mux_1314_i27_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[26]), 
         .D(n224[26]), .Z(n3181[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i27_3_lut_4_lut.init = 16'hf780;
    LUT4 reduce_or_459_i1_3_lut (.A(busy), .B(n1286[13]), .C(n1286[20]), 
         .Z(n1397)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam reduce_or_459_i1_3_lut.init = 16'hdcdc;
    FD1P3IX esc_data_i0_i3 (.D(n9241[3]), .SP(n12098), .CD(n14425), .CK(debug_c_c), 
            .Q(esc_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i3.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i5 (.D(n9241[5]), .SP(n12098), .CD(n14425), .CK(debug_c_c), 
            .Q(esc_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i5.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i6 (.D(n9241[6]), .SP(n12098), .CD(n14425), .CK(debug_c_c), 
            .Q(esc_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i6.GSR = "ENABLED";
    FD1P3IX esc_data_i0_i7 (.D(n9241[7]), .SP(n12098), .CD(n14425), .CK(debug_c_c), 
            .Q(esc_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i7.GSR = "ENABLED";
    LUT4 mux_1314_i26_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[25]), 
         .D(n224[25]), .Z(n3181[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i26_3_lut_4_lut.init = 16'hf780;
    FD1P3AX select__i1 (.D(n29730), .SP(n12788), .CK(debug_c_c), .Q(\select[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i1.GSR = "ENABLED";
    LUT4 i24473_then_3_lut (.A(\buffer[0] [7]), .B(\buffer[2] [7]), .C(\sendcount[1] ), 
         .Z(n32523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24473_then_3_lut.init = 16'hcaca;
    LUT4 i24473_else_3_lut (.A(\buffer[3] [7]), .B(\buffer[1] [7]), .C(\sendcount[1] ), 
         .Z(n32522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24473_else_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(esc_data[1]), .B(esc_data[3]), .C(esc_data[4]), 
         .D(esc_data[2]), .Z(n35)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut.init = 16'h5f4c;
    LUT4 i4_4_lut (.A(rx_data[2]), .B(n30114), .C(rx_data[5]), .D(n6_c), 
         .Z(n11639)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i4_4_lut.init = 16'h0800;
    LUT4 i498_2_lut (.A(n1286[3]), .B(n1286[4]), .Z(n1687)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i498_2_lut.init = 16'heeee;
    LUT4 i2_4_lut (.A(escape), .B(n13_c), .C(debug_c_7), .D(n11539), 
         .Z(n30114)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i2_4_lut.init = 16'h1000;
    LUT4 i1_2_lut (.A(n1286[3]), .B(rx_data[0]), .Z(n6_c)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i24476_then_3_lut (.A(\buffer[0] [6]), .B(\buffer[2] [6]), .C(\sendcount[1] ), 
         .Z(n32526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24476_then_3_lut.init = 16'hcaca;
    LUT4 i24476_else_3_lut (.A(\buffer[3] [6]), .B(\buffer[1] [6]), .C(\sendcount[1] ), 
         .Z(n32525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24476_else_3_lut.init = 16'hcaca;
    LUT4 equal_143_i13_2_lut (.A(rx_data[6]), .B(rx_data[7]), .Z(n13_c)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(139[12:17])
    defparam equal_143_i13_2_lut.init = 16'heeee;
    LUT4 i24479_then_3_lut (.A(\buffer[0] [5]), .B(\buffer[2] [5]), .C(\sendcount[1] ), 
         .Z(n32529)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24479_then_3_lut.init = 16'hcaca;
    LUT4 i24780_3_lut (.A(debug_c_7), .B(n29974), .C(n1286[3]), .Z(n30109)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i24780_3_lut.init = 16'h2020;
    LUT4 i24479_else_3_lut (.A(\buffer[3] [5]), .B(\buffer[1] [5]), .C(\sendcount[1] ), 
         .Z(n32528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24479_else_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut (.A(n30619), .B(n31474), .C(rx_data[0]), .D(escape), 
         .Z(n29974)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut.init = 16'h0040;
    LUT4 i4986_3_lut (.A(debug_c_7), .B(n1286[3]), .C(n1286[2]), .Z(n10751)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4986_3_lut.init = 16'h5454;
    LUT4 i1_4_lut_adj_68 (.A(n1286[4]), .B(debug_c_7), .C(n1286[2]), .D(n30106), 
         .Z(n29412)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_68.init = 16'heeea;
    LUT4 i1_4_lut_adj_69 (.A(n15_c), .B(n1286[3]), .C(n1318), .D(n30714), 
         .Z(n30106)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (C+!(D))+!B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_69.init = 16'h50dc;
    LUT4 i24482_then_3_lut (.A(\buffer[0] [4]), .B(\buffer[2] [4]), .C(\sendcount[1] ), 
         .Z(n32532)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24482_then_3_lut.init = 16'hcaca;
    LUT4 i24355_3_lut (.A(n11477), .B(escape), .C(n15_c), .Z(n30714)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24355_3_lut.init = 16'hecec;
    LUT4 i2_4_lut_adj_70 (.A(n29621), .B(rx_data[4]), .C(rx_data[1]), 
         .D(rx_data[3]), .Z(n11477)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(150[12:17])
    defparam i2_4_lut_adj_70.init = 16'hbfff;
    LUT4 i3_4_lut_adj_71 (.A(rx_data[4]), .B(rx_data[3]), .C(rx_data[1]), 
         .D(n29621), .Z(n15_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(150[12:17])
    defparam i3_4_lut_adj_71.init = 16'hfffe;
    LUT4 i13994_2_lut (.A(bufcount[1]), .B(n1318), .Z(n14082)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i13994_2_lut.init = 16'h2222;
    LUT4 i24482_else_3_lut (.A(\buffer[3] [4]), .B(\buffer[1] [4]), .C(\sendcount[1] ), 
         .Z(n32531)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24482_else_3_lut.init = 16'hcaca;
    LUT4 mux_1314_i25_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[24]), 
         .D(n224[24]), .Z(n3181[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i25_3_lut_4_lut.init = 16'hf780;
    LUT4 i14770_3_lut_rep_327 (.A(n2497), .B(n32444), .C(n1286[18]), .Z(n32421)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i14770_3_lut_rep_327.init = 16'hc8c8;
    FD1P3AX select__i2 (.D(n29727), .SP(n12788), .CK(debug_c_c), .Q(\select[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i2.GSR = "ENABLED";
    FD1P3AX select__i4 (.D(n29726), .SP(n12788), .CK(debug_c_c), .Q(\select[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i4.GSR = "ENABLED";
    FD1P3AX select__i7 (.D(n30279), .SP(n12788), .CK(debug_c_c), .Q(\select[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam select__i7.GSR = "ENABLED";
    LUT4 i24648_2_lut_3_lut (.A(n2497), .B(n32444), .C(n1286[18]), .Z(n14122)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i24648_2_lut_3_lut.init = 16'h0808;
    LUT4 i14436_4_lut (.A(sendcount[2]), .B(n32380), .C(n9_c), .D(n32464), 
         .Z(n18[2])) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+!((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i14436_4_lut.init = 16'h1323;
    LUT4 i25222_then_3_lut (.A(\buffer[0] [0]), .B(\buffer[2] [0]), .C(\sendcount[1] ), 
         .Z(n32535)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25222_then_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_72 (.A(n13_c), .B(rx_data[5]), .C(rx_data[2]), .D(rx_data[0]), 
         .Z(n29621)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(150[12:17])
    defparam i2_4_lut_adj_72.init = 16'hfeff;
    LUT4 i25222_else_3_lut (.A(\buffer[3] [0]), .B(\buffer[1] [0]), .C(\sendcount[1] ), 
         .Z(n32534)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i25222_else_3_lut.init = 16'hcaca;
    FD1P3AX sendcount__i2 (.D(n18[2]), .SP(n32407), .CK(debug_c_c), .Q(sendcount[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i2.GSR = "ENABLED";
    FD1P3IX sendcount__i1 (.D(n19[1]), .SP(n32407), .CD(n32380), .CK(debug_c_c), 
            .Q(\sendcount[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i1.GSR = "ENABLED";
    LUT4 n30389_bdd_4_lut (.A(sendcount[3]), .B(sendcount[2]), .C(sendcount[0]), 
         .D(\sendcount[1] ), .Z(n31398)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam n30389_bdd_4_lut.init = 16'h4001;
    LUT4 n32270_bdd_3_lut_4_lut (.A(sendcount[2]), .B(n32476), .C(n32536), 
         .D(n32270), .Z(n32271)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam n32270_bdd_3_lut_4_lut.init = 16'hf960;
    LUT4 mux_429_Mux_7_i7_4_lut_4_lut (.A(n32515), .B(n32461), .C(n4_adj_28), 
         .D(n32524), .Z(n9241[7])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_7_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i1_4_lut_adj_73 (.A(n32463), .B(debug_c_7), .C(n11639), .D(n8), 
         .Z(n29464)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_73.init = 16'hdc50;
    LUT4 mux_1314_i24_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[23]), 
         .D(n224[23]), .Z(n3181[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i23_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[22]), 
         .D(n224[22]), .Z(n3181[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i22_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[21]), 
         .D(n224[21]), .Z(n3181[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 i13969_2_lut (.A(bufcount[0]), .B(n1318), .Z(n13423)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i13969_2_lut.init = 16'h2222;
    LUT4 i24485_then_3_lut (.A(\buffer[0] [3]), .B(\buffer[2] [3]), .C(\sendcount[1] ), 
         .Z(n32538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24485_then_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut (.A(n15_c), .B(n1286[1]), .C(n1318), .Z(n8)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_3_lut.init = 16'hecec;
    LUT4 mux_429_Mux_6_i7_4_lut_4_lut (.A(n32515), .B(n32461), .C(n4_adj_29), 
         .D(n32527), .Z(n9241[6])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_6_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_5_i7_4_lut_4_lut (.A(n32515), .B(n32461), .C(n4_adj_30), 
         .D(n32530), .Z(n9241[5])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_5_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 mux_429_Mux_3_i7_4_lut_4_lut (.A(n32515), .B(n32461), .C(n4_adj_31), 
         .D(n32539), .Z(n9241[3])) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam mux_429_Mux_3_i7_4_lut_4_lut.init = 16'hdc10;
    LUT4 i24485_else_3_lut (.A(\buffer[3] [3]), .B(\buffer[1] [3]), .C(\sendcount[1] ), 
         .Z(n32537)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24485_else_3_lut.init = 16'hcaca;
    LUT4 mux_1314_i21_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[20]), 
         .D(n224[20]), .Z(n3181[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 i24488_then_3_lut (.A(\buffer[0] [2]), .B(\buffer[2] [2]), .C(\sendcount[1] ), 
         .Z(n32541)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24488_then_3_lut.init = 16'hcaca;
    LUT4 mux_1314_i20_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[19]), 
         .D(n224[19]), .Z(n3181[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 i24488_else_3_lut (.A(\buffer[3] [2]), .B(\buffer[1] [2]), .C(\sendcount[1] ), 
         .Z(n32540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24488_else_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(n1286[4]), .B(n32469), .C(bufcount[0]), 
         .D(n32445), .Z(n28389)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'hd222;
    LUT4 mux_1314_i19_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[18]), 
         .D(n224[18]), .Z(n3181[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 i24491_then_3_lut (.A(\buffer[0] [1]), .B(\buffer[2] [1]), .C(\sendcount[1] ), 
         .Z(n32544)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24491_then_3_lut.init = 16'hcaca;
    LUT4 mux_1314_i18_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[17]), 
         .D(n224[17]), .Z(n3181[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32468), .B(bufcount[3]), .C(\buffer[0] [7]), 
         .D(n11639), .Z(n30166)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0e00;
    LUT4 mux_1314_i17_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[16]), 
         .D(n224[16]), .Z(n3181[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i16_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[15]), 
         .D(n224[15]), .Z(n3181[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 i2992_2_lut_rep_370 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n32464)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2992_2_lut_rep_370.init = 16'h8888;
    LUT4 i2891_2_lut_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(sendcount[2]), 
         .Z(n8679)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2891_2_lut_3_lut.init = 16'h8080;
    LUT4 i24491_else_3_lut (.A(\buffer[3] [1]), .B(\buffer[1] [1]), .C(\sendcount[1] ), 
         .Z(n32543)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24491_else_3_lut.init = 16'hcaca;
    LUT4 mux_1314_i15_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[14]), 
         .D(n224[14]), .Z(n3181[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 i8325_then_4_lut (.A(bufcount[3]), .B(n1318), .C(n1286[3]), .D(n1286[4]), 
         .Z(n32547)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i8325_then_4_lut.init = 16'haaa2;
    LUT4 i8325_else_4_lut (.A(bufcount[3]), .B(n1318), .C(n1286[3]), .D(n1286[4]), 
         .Z(n32546)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i8325_else_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_adj_74 (.A(register_addr[1]), .B(\steps_reg[4] ), .Z(n15)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_74.init = 16'h8888;
    LUT4 mux_1314_i14_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[13]), 
         .D(n224[13]), .Z(n3181[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i13_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[12]), 
         .D(n224[12]), .Z(n3181[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 n33741_bdd_4_lut (.A(n33741), .B(n1286[4]), .C(n33743), .D(bufcount[2]), 
         .Z(n34314)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n33741_bdd_4_lut.init = 16'heef0;
    LUT4 mux_1314_i12_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[11]), 
         .D(n224[11]), .Z(n3181[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_75 (.A(n9), .B(n8204[0]), .C(n32444), .D(n1304), 
         .Z(n14425)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_75.init = 16'h8000;
    LUT4 mux_1384_i13_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[12]), 
         .D(n224_adj_42[12]), .Z(n3451[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i11_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[10]), 
         .D(n224[10]), .Z(n3181[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i10_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[9]), 
         .D(n224[9]), .Z(n3181[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_76 (.A(register_addr[1]), .B(\steps_reg[7] ), .Z(n13)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_76.init = 16'h8888;
    LUT4 mux_429_Mux_3_i4_3_lut (.A(\buffer[4] [3]), .B(\buffer[5] [3]), 
         .C(sendcount[0]), .Z(n4_adj_31)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_3_i4_3_lut.init = 16'hacac;
    LUT4 mux_1384_i12_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[11]), 
         .D(n224_adj_42[11]), .Z(n3451[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i11_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[10]), 
         .D(n224_adj_42[10]), .Z(n3451[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i9_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[8]), 
         .D(n224[8]), .Z(n3181[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i10_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[9]), 
         .D(n224_adj_42[9]), .Z(n3451[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i9_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[8]), 
         .D(n224_adj_42[8]), .Z(n3451[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i8_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[7]), 
         .D(n224_adj_42[7]), .Z(n3451[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i7_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[6]), 
         .D(n224_adj_42[6]), .Z(n3451[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_429_Mux_5_i4_3_lut (.A(\buffer[4] [5]), .B(\buffer[5] [5]), 
         .C(sendcount[0]), .Z(n4_adj_30)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_5_i4_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_adj_77 (.A(register_addr[1]), .B(\steps_reg[3] ), .Z(n15_adj_33)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_77.init = 16'h8888;
    LUT4 i2838_2_lut_3_lut_4_lut_4_lut (.A(bufcount[1]), .B(n32445), .C(n32462), 
         .D(bufcount[0]), .Z(n1682[1])) /* synthesis lut_function=(A (B (C+!(D)))+!A !((C+!(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i2838_2_lut_3_lut_4_lut_4_lut.init = 16'h8488;
    FD1P3AX rw_498 (.D(n1286[10]), .SP(n2539), .CK(debug_c_c), .Q(rw));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498.GSR = "ENABLED";
    LUT4 mux_1384_i6_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[5]), 
         .D(n224_adj_42[5]), .Z(n3451[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 i2787_2_lut_rep_374 (.A(bufcount[1]), .B(bufcount[2]), .Z(n32468)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2787_2_lut_rep_374.init = 16'heeee;
    LUT4 mux_1384_i5_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[4]), 
         .D(n224_adj_42[4]), .Z(n3451[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i5_3_lut_4_lut.init = 16'hf780;
    FD1S3AX escape_501 (.D(n9337), .CK(debug_c_c), .Q(escape));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam escape_501.GSR = "ENABLED";
    LUT4 mux_1314_i8_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[7]), 
         .D(n224[7]), .Z(n3181[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_78 (.A(register_addr[1]), .B(\steps_reg[5] ), .Z(n14)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_78.init = 16'h8888;
    LUT4 mux_1384_i4_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[3]), 
         .D(n224_adj_42[3]), .Z(n3451[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut (.A(n1286[3]), .B(n30754), .C(\buffer[2] [4]), 
         .Z(n30175)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_79 (.A(n1286[3]), .B(n30754), .C(\buffer[2] [3]), 
         .Z(n30179)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_79.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_80 (.A(n1286[3]), .B(n30754), .C(\buffer[2] [2]), 
         .Z(n30184)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_80.init = 16'h8080;
    LUT4 i2424_2_lut_rep_369_3_lut (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[3]), 
         .Z(n32463)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2424_2_lut_rep_369_3_lut.init = 16'hfefe;
    LUT4 mux_1314_i7_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[6]), 
         .D(n224[6]), .Z(n3181[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_adj_81 (.A(n1286[3]), .B(n30754), .C(\buffer[2] [1]), 
         .Z(n30177)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_81.init = 16'h8080;
    LUT4 mux_429_Mux_6_i4_3_lut (.A(\buffer[4] [6]), .B(\buffer[5] [6]), 
         .C(sendcount[0]), .Z(n4_adj_29)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_6_i4_3_lut.init = 16'hacac;
    LUT4 mux_1384_i3_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[2]), 
         .D(n224_adj_42[2]), .Z(n3451[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_adj_82 (.A(n1286[3]), .B(n30754), .C(\buffer[2] [0]), 
         .Z(n30183)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_82.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_83 (.A(n1286[3]), .B(n30754), .C(n1286[13]), 
         .Z(n14_adj_43)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_83.init = 16'hf8f8;
    LUT4 mux_1384_i2_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[1]), 
         .D(n224_adj_42[1]), .Z(n3451[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_adj_84 (.A(n1286[3]), .B(n30754), .C(\buffer[2] [5]), 
         .Z(n30182)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_84.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_85 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n30487)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_85.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_86 (.A(n1286[3]), .B(n30754), .C(\buffer[2] [6]), 
         .Z(n30185)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_86.init = 16'h8080;
    LUT4 mux_1314_i6_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[5]), 
         .D(n224[5]), .Z(n3181[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_adj_87 (.A(bufcount[1]), .B(bufcount[2]), .C(bufcount[0]), 
         .Z(n30488)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_87.init = 16'hbfbf;
    LUT4 mux_1314_i5_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[4]), 
         .D(n224[4]), .Z(n3181[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i32_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[31]), 
         .D(n224_adj_42[31]), .Z(n3451[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i32_3_lut_4_lut.init = 16'hf780;
    LUT4 i14662_3_lut_rep_375 (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .Z(n32469)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i14662_3_lut_rep_375.init = 16'hecec;
    LUT4 i1_2_lut_3_lut_adj_88 (.A(n1286[3]), .B(n30754), .C(\buffer[2] [7]), 
         .Z(n30186)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_88.init = 16'h8080;
    LUT4 i2_2_lut_rep_368_4_lut (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1286[4]), .Z(n32462)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+!(D))) */ ;
    defparam i2_2_lut_rep_368_4_lut.init = 16'hecff;
    LUT4 i1_2_lut_4_lut (.A(bufcount[1]), .B(bufcount[3]), .C(bufcount[2]), 
         .D(n1286[4]), .Z(n7)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hec00;
    LUT4 i854_2_lut_rep_376 (.A(escape), .B(debug_c_7), .Z(n32470)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i854_2_lut_rep_376.init = 16'hbbbb;
    LUT4 mux_1384_i31_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[30]), 
         .D(n224_adj_42[30]), .Z(n3451[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i31_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_3_lut_rep_351_4_lut (.A(escape), .B(debug_c_7), .C(n30754), 
         .D(n1286[4]), .Z(n32445)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(125[8] 167[12])
    defparam i2_3_lut_rep_351_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut_3_lut_adj_89 (.A(n1286[3]), .B(n30754), .C(\buffer[3] [0]), 
         .Z(n30187)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_89.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_90 (.A(n1286[3]), .B(n30754), .C(\buffer[3] [1]), 
         .Z(n30188)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_90.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_91 (.A(n1286[3]), .B(n30754), .C(\buffer[3] [2]), 
         .Z(n30189)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_91.init = 16'h8080;
    LUT4 mux_429_Mux_7_i4_3_lut (.A(\buffer[4] [7]), .B(\buffer[5] [7]), 
         .C(sendcount[0]), .Z(n4_adj_28)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_7_i4_3_lut.init = 16'hacac;
    LUT4 mux_1314_i4_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[3]), 
         .D(n224[3]), .Z(n3181[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_adj_92 (.A(n1286[3]), .B(n30754), .C(\buffer[3] [3]), 
         .Z(n30193)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_92.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_93 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n30512)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_93.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_94 (.A(n1286[3]), .B(n30754), .C(\buffer[3] [4]), 
         .Z(n30178)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_94.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_95 (.A(bufcount[2]), .B(bufcount[1]), .C(bufcount[0]), 
         .Z(n30511)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(176[12:28])
    defparam i1_2_lut_3_lut_adj_95.init = 16'hbfbf;
    LUT4 i1_2_lut_3_lut_adj_96 (.A(n1286[3]), .B(n30754), .C(\buffer[3] [5]), 
         .Z(n30192)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_96.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_97 (.A(n1286[3]), .B(n30754), .C(\buffer[3] [6]), 
         .Z(n30194)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_97.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_98 (.A(n1286[3]), .B(n30754), .C(\buffer[3] [7]), 
         .Z(n30191)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_98.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_99 (.A(n1286[3]), .B(n30754), .C(\buffer[4] [0]), 
         .Z(n30190)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_99.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_100 (.A(n1286[3]), .B(n30754), .C(\buffer[4] [1]), 
         .Z(n30181)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_100.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_101 (.A(n1286[3]), .B(n30754), .C(\buffer[4] [2]), 
         .Z(n30195)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_101.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_102 (.A(n1286[3]), .B(n30754), .C(\buffer[4] [3]), 
         .Z(n30196)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_102.init = 16'h8080;
    LUT4 mux_1314_i3_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[2]), 
         .D(n224[2]), .Z(n3181[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_4_lut_adj_103 (.A(databus[19]), .B(n5_c), .C(n1286[13]), .D(n30196), 
         .Z(n28336)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_103.init = 16'hffec;
    LUT4 i1_2_lut_3_lut_adj_104 (.A(n1286[3]), .B(n30754), .C(\buffer[4] [4]), 
         .Z(n30198)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_104.init = 16'h8080;
    LUT4 mux_1384_i30_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[29]), 
         .D(n224_adj_42[29]), .Z(n3451[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i30_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_adj_105 (.A(n1286[3]), .B(n30754), .C(\buffer[4] [5]), 
         .Z(n30180)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_105.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_106 (.A(n1286[3]), .B(n30754), .C(\buffer[4] [6]), 
         .Z(n30197)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_106.init = 16'h8080;
    LUT4 mux_1314_i2_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[1]), 
         .D(n224[1]), .Z(n3181[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_512_i1_3_lut (.A(n2497), .B(esc_data[0]), .C(n1286[18]), 
         .Z(n2028[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_512_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_107 (.A(n1286[3]), .B(n30754), .C(\buffer[4] [7]), 
         .Z(n30201)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_107.init = 16'h8080;
    LUT4 i1_2_lut_rep_381 (.A(n1304), .B(sendcount[4]), .Z(n32475)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_381.init = 16'h2222;
    LUT4 select_1742_Select_35_i5_4_lut (.A(\buffer[4] [3]), .B(n1286[4]), 
         .C(rx_data[3]), .D(n30487), .Z(n5_c)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_35_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_108 (.A(n1286[3]), .B(n30754), .C(\buffer[5] [0]), 
         .Z(n30200)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_108.init = 16'h8080;
    LUT4 i1_2_lut_adj_109 (.A(sendcount[0]), .B(sendcount[3]), .Z(n4)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_109.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_110 (.A(n1286[3]), .B(n30754), .C(\buffer[5] [1]), 
         .Z(n30176)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_110.init = 16'h8080;
    FD1P3AX sendcount__i3 (.D(n28153), .SP(n32407), .CK(debug_c_c), .Q(sendcount[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i3.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_111 (.A(n1286[3]), .B(n30754), .C(\buffer[5] [2]), 
         .Z(n30202)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_111.init = 16'h8080;
    FD1P3AX sendcount__i4 (.D(n17), .SP(n32407), .CK(debug_c_c), .Q(sendcount[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam sendcount__i4.GSR = "ENABLED";
    LUT4 expansion5_c_bdd_2_lut_24899_3_lut (.A(n1304), .B(sendcount[4]), 
         .C(n31398), .Z(n31399)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam expansion5_c_bdd_2_lut_24899_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_112 (.A(n1286[3]), .B(n30754), .C(\buffer[5] [3]), 
         .Z(n30203)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_112.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_113 (.A(n1286[3]), .B(n30754), .C(\buffer[5] [4]), 
         .Z(n30204)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_113.init = 16'h8080;
    LUT4 i13875_2_lut_rep_382 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n32476)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13875_2_lut_rep_382.init = 16'heeee;
    LUT4 i1_2_lut_rep_367_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(sendcount[2]), 
         .Z(n32461)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam i1_2_lut_rep_367_3_lut.init = 16'h1e1e;
    LUT4 i1_2_lut_3_lut_adj_114 (.A(n1286[3]), .B(n30754), .C(\buffer[5] [5]), 
         .Z(n30206)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_114.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_115 (.A(n1286[3]), .B(n30754), .C(\buffer[5] [6]), 
         .Z(n30199)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_115.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_116 (.A(n1286[3]), .B(n30754), .C(\buffer[5] [7]), 
         .Z(n30205)) /* synthesis lut_function=(A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_116.init = 16'h8080;
    LUT4 mux_1384_i29_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[28]), 
         .D(n224_adj_42[28]), .Z(n3451[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i29_3_lut_4_lut.init = 16'hf780;
    LUT4 i4_2_lut_rep_384 (.A(n1304), .B(n1286[15]), .Z(n32478)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_2_lut_rep_384.init = 16'heeee;
    LUT4 i2_4_lut_adj_117 (.A(databus[20]), .B(n5_adj_50), .C(n1286[13]), 
         .D(n30198), .Z(n28343)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_117.init = 16'hffec;
    LUT4 i1_2_lut_3_lut_adj_118 (.A(n1304), .B(n1286[15]), .C(n1286[12]), 
         .Z(n30537)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_118.init = 16'hfefe;
    LUT4 i51_4_lut (.A(esc_data[2]), .B(esc_data[3]), .C(esc_data[4]), 
         .D(esc_data[1]), .Z(n55)) /* synthesis lut_function=(A (B)+!A !(B+!(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i51_4_lut.init = 16'h9998;
    LUT4 select_1742_Select_36_i5_4_lut (.A(\buffer[4] [4]), .B(n1286[4]), 
         .C(rx_data[4]), .D(n30487), .Z(n5_adj_50)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_36_i5_4_lut.init = 16'h88c0;
    LUT4 mux_1384_i20_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[19]), 
         .D(n224_adj_42[19]), .Z(n3451[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i19_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[18]), 
         .D(n224_adj_42[18]), .Z(n3451[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i28_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[27]), 
         .D(n224_adj_42[27]), .Z(n3451[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i28_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_119 (.A(n1286[4]), .B(\buffer[0] [6]), .C(n11_adj_10), 
         .D(n14_adj_43), .Z(n29260)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_119.init = 16'heca0;
    LUT4 i13873_2_lut (.A(sendcount[3]), .B(sendcount[0]), .Z(n8204[0])) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i13873_2_lut.init = 16'hdddd;
    LUT4 n11281_bdd_2_lut (.A(sendcount[0]), .B(sendcount[3]), .Z(n32266)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam n11281_bdd_2_lut.init = 16'hbbbb;
    LUT4 i884_2_lut (.A(n1286[5]), .B(n32444), .Z(n2541)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(88[5] 327[8])
    defparam i884_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_388 (.A(n1286[3]), .B(n1286[19]), .Z(n32482)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_388.init = 16'heeee;
    LUT4 i1_2_lut_rep_389 (.A(n1286[11]), .B(n1286[9]), .Z(n32483)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_389.init = 16'heeee;
    LUT4 i3_2_lut_3_lut_4_lut (.A(n1286[11]), .B(n1286[9]), .C(n1286[19]), 
         .D(n1286[3]), .Z(n9_adj_53)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_1384_i27_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[26]), 
         .D(n224_adj_42[26]), .Z(n3451[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i27_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i26_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[25]), 
         .D(n224_adj_42[25]), .Z(n3451[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i26_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_3_lut_rep_390 (.A(n1286[13]), .B(n1286[7]), .C(n1286[5]), 
         .Z(n32484)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_3_lut_rep_390.init = 16'hfefe;
    LUT4 mux_1314_i28_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[27]), 
         .D(n224[27]), .Z(n3181[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i28_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_2_lut_4_lut (.A(n1286[13]), .B(n1286[7]), .C(n1286[5]), .D(n1286[17]), 
         .Z(n8_adj_57)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_2_lut_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_120 (.A(databus[21]), .B(n5_adj_58), .C(n1286[13]), 
         .D(n30180), .Z(n28341)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_120.init = 16'hffec;
    LUT4 i2_4_lut_adj_121 (.A(\buffer[0] [2]), .B(\buffer[0] [0]), .C(n30278), 
         .D(\buffer[0] [1]), .Z(n29730)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i2_4_lut_adj_121.init = 16'h0040;
    LUT4 i1_4_lut_adj_122 (.A(\buffer[0] [3]), .B(n18427), .C(n6_adj_59), 
         .D(\buffer[0] [4]), .Z(n30278)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_122.init = 16'h0004;
    LUT4 i2_2_lut (.A(\buffer[0] [5]), .B(\buffer[0] [6]), .Z(n6_adj_59)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(227[9:31])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 mux_1384_i25_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[24]), 
         .D(n224_adj_42[24]), .Z(n3451[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i25_3_lut_4_lut.init = 16'hf780;
    FD1P3AX send_491 (.D(n11238), .SP(n28369), .CK(debug_c_c), .Q(send));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam send_491.GSR = "ENABLED";
    PFUMX i25259 (.BLUT(n32516), .ALUT(n32517), .C0(sendcount[3]), .Z(n9));
    LUT4 i2_4_lut_adj_123 (.A(databus[1]), .B(n5_adj_61), .C(n1286[13]), 
         .D(n30177), .Z(n28235)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_123.init = 16'hffec;
    LUT4 mux_512_i5_3_lut (.A(n2497), .B(esc_data[4]), .C(n1286[18]), 
         .Z(n2028[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_512_i5_3_lut.init = 16'hcaca;
    LUT4 select_1742_Select_17_i5_4_lut (.A(\buffer[2] [1]), .B(n1286[4]), 
         .C(rx_data[1]), .D(n30512), .Z(n5_adj_61)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_17_i5_4_lut.init = 16'h88c0;
    LUT4 mux_1384_i24_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[23]), 
         .D(n224_adj_42[23]), .Z(n3451[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 select_1742_Select_37_i5_4_lut (.A(\buffer[4] [5]), .B(n1286[4]), 
         .C(rx_data[5]), .D(n30487), .Z(n5_adj_58)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_37_i5_4_lut.init = 16'h88c0;
    LUT4 mux_1384_i23_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[22]), 
         .D(n224_adj_42[22]), .Z(n3451[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 i4912_3_lut (.A(busy), .B(n1286[17]), .C(n1286[16]), .Z(n10675)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4912_3_lut.init = 16'ha8a8;
    LUT4 i1_4_lut_then_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(\sendcount[1] ), 
         .D(sendcount[2]), .Z(n32517)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i1_4_lut_then_4_lut.init = 16'h0001;
    LUT4 i2_4_lut_adj_124 (.A(n30278), .B(\buffer[0] [0]), .C(\buffer[0] [2]), 
         .D(\buffer[0] [1]), .Z(n30279)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_4_lut_adj_124.init = 16'h8000;
    LUT4 mux_1384_i18_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[17]), 
         .D(n224_adj_42[17]), .Z(n3451[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 i5_4_lut (.A(esc_data[0]), .B(n10), .C(n30705), .D(n30), .Z(n2497)) /* synthesis lut_function=(A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i5_4_lut.init = 16'h8808;
    LUT4 sendcount_4__bdd_3_lut_25128 (.A(sendcount[4]), .B(n31947), .C(sendcount[3]), 
         .Z(n31948)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam sendcount_4__bdd_3_lut_25128.init = 16'hcaca;
    LUT4 i2_4_lut_adj_125 (.A(databus[22]), .B(n5_adj_65), .C(n1286[13]), 
         .D(n30197), .Z(n28338)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_125.init = 16'hffec;
    LUT4 mux_1384_i22_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[21]), 
         .D(n224_adj_42[21]), .Z(n3451[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 i4_4_lut_adj_126 (.A(n1286[15]), .B(esc_data[6]), .C(esc_data[5]), 
         .D(esc_data[7]), .Z(n10)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut_adj_126.init = 16'h0002;
    LUT4 select_1742_Select_38_i5_4_lut (.A(\buffer[4] [6]), .B(n1286[4]), 
         .C(rx_data[6]), .D(n30487), .Z(n5_adj_65)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_38_i5_4_lut.init = 16'h88c0;
    LUT4 sendcount_4__bdd_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(sendcount[2]), 
         .D(\sendcount[1] ), .Z(n31947)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;
    defparam sendcount_4__bdd_4_lut.init = 16'h6aaa;
    LUT4 mux_1384_i21_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[20]), 
         .D(n224_adj_42[20]), .Z(n3451[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1384_i17_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[16]), 
         .D(n224_adj_42[16]), .Z(n3451[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i17_3_lut_4_lut.init = 16'hf780;
    FD1P3IX tx_data_i0_i2 (.D(esc_data[2]), .SP(n32421), .CD(n14122), 
            .CK(debug_c_c), .Q(tx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i2.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i5 (.D(esc_data[5]), .SP(n32421), .CD(n14122), 
            .CK(debug_c_c), .Q(tx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i5.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i6 (.D(esc_data[6]), .SP(n32421), .CD(n14122), 
            .CK(debug_c_c), .Q(tx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i6.GSR = "ENABLED";
    FD1P3IX tx_data_i0_i7 (.D(esc_data[7]), .SP(n32421), .CD(n14122), 
            .CK(debug_c_c), .Q(tx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam tx_data_i0_i7.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_127 (.A(n1286[4]), .B(\buffer[0] [5]), .C(n11_adj_11), 
         .D(n14_adj_43), .Z(n29262)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_127.init = 16'heca0;
    LUT4 i2_4_lut_adj_128 (.A(databus[23]), .B(n5_adj_69), .C(n1286[13]), 
         .D(n30201), .Z(n28305)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_128.init = 16'hffec;
    LUT4 i24347_4_lut (.A(esc_data[4]), .B(esc_data[1]), .C(esc_data[3]), 
         .D(esc_data[2]), .Z(n30705)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24347_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_129 (.A(esc_data[1]), .B(esc_data[2]), .C(esc_data[4]), 
         .D(esc_data[3]), .Z(n30)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_129.init = 16'h2080;
    LUT4 mux_512_i4_3_lut (.A(n2497), .B(esc_data[3]), .C(n1286[18]), 
         .Z(n2028[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_512_i4_3_lut.init = 16'hcaca;
    LUT4 mux_512_i2_3_lut (.A(n2497), .B(esc_data[1]), .C(n1286[18]), 
         .Z(n2028[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam mux_512_i2_3_lut.init = 16'hcaca;
    LUT4 select_1742_Select_39_i5_4_lut (.A(\buffer[4] [7]), .B(n1286[4]), 
         .C(rx_data[7]), .D(n30487), .Z(n5_adj_69)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_39_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_130 (.A(databus[24]), .B(n5_adj_70), .C(n1286[13]), 
         .D(n30200), .Z(n28358)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_130.init = 16'hffec;
    LUT4 i1_4_lut_adj_131 (.A(n1286[4]), .B(\buffer[0] [4]), .C(n11_adj_12), 
         .D(n14_adj_43), .Z(n29266)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_131.init = 16'heca0;
    LUT4 select_1742_Select_40_i5_4_lut (.A(\buffer[5] [0]), .B(n1286[4]), 
         .C(rx_data[0]), .D(n30488), .Z(n5_adj_70)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_40_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut_adj_132 (.A(n1286[4]), .B(\buffer[0] [3]), .C(n11_adj_13), 
         .D(n14_adj_43), .Z(n29326)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_132.init = 16'heca0;
    FD1P3AX databus_out_i0_i31 (.D(\buffer[5] [7]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i31.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i30 (.D(\buffer[5] [6]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i30.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i29 (.D(\buffer[5] [5]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i29.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i28 (.D(\buffer[5] [4]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i28.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i27 (.D(\buffer[5] [3]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i27.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i26 (.D(\buffer[5] [2]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i26.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i25 (.D(\buffer[5] [1]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i25.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i24 (.D(\buffer[5] [0]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i24.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i23 (.D(\buffer[4] [7]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i23.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i22 (.D(\buffer[4] [6]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i22.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i21 (.D(\buffer[4] [5]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i21.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i20 (.D(\buffer[4] [4]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i20.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i19 (.D(\buffer[4] [3]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i19.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i18 (.D(\buffer[4] [2]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i18.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i17 (.D(\buffer[4] [1]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i17.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i16 (.D(\buffer[4] [0]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i16.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i15 (.D(\buffer[3] [7]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i15.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_133 (.A(databus[25]), .B(n5_adj_71), .C(n1286[13]), 
         .D(n30176), .Z(n28370)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_133.init = 16'hffec;
    FD1P3AX databus_out_i0_i14 (.D(\buffer[3] [6]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i14.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i13 (.D(\buffer[3] [5]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i13.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i12 (.D(\buffer[3] [4]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i12.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i11 (.D(\buffer[3] [3]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i11.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i10 (.D(\buffer[3] [2]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i10.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i9 (.D(\buffer[3] [1]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i9.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i8 (.D(\buffer[3] [0]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i8.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i7 (.D(\buffer[2] [7]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i7.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i6 (.D(\buffer[2] [6]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i6.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i5 (.D(\buffer[2] [5]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i5.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i4 (.D(\buffer[2] [4]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i4.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i3 (.D(\buffer[2] [3]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i3.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i2 (.D(\buffer[2] [2]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i2.GSR = "ENABLED";
    FD1P3AX databus_out_i0_i1 (.D(\buffer[2] [1]), .SP(n2541), .CK(debug_c_c), 
            .Q(databus_out[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam databus_out_i0_i1.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i4 (.D(n4846[4]), .SP(n12098), .CK(debug_c_c), 
            .Q(esc_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i4.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i2 (.D(n4846[2]), .SP(n12098), .CK(debug_c_c), 
            .Q(esc_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i2.GSR = "ENABLED";
    FD1P3AX esc_data_i0_i1 (.D(n4846[1]), .SP(n12098), .CK(debug_c_c), 
            .Q(esc_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam esc_data_i0_i1.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_134 (.A(n1286[4]), .B(\buffer[0] [2]), .C(n11_adj_14), 
         .D(n14_adj_43), .Z(n29198)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_134.init = 16'heca0;
    LUT4 select_1742_Select_41_i5_4_lut (.A(\buffer[5] [1]), .B(n1286[4]), 
         .C(rx_data[1]), .D(n30488), .Z(n5_adj_71)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_41_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut_adj_135 (.A(n1286[4]), .B(\buffer[0] [1]), .C(n11_adj_15), 
         .D(n14_adj_43), .Z(n29186)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_135.init = 16'heca0;
    LUT4 i3680_3_lut (.A(n1286[16]), .B(n2497), .C(busy), .Z(n9441)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3680_3_lut.init = 16'hcece;
    LUT4 i1_4_lut_else_4_lut (.A(sendcount[4]), .B(sendcount[0]), .C(\sendcount[1] ), 
         .D(sendcount[2]), .Z(n32516)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam i1_4_lut_else_4_lut.init = 16'h4001;
    LUT4 n30754_bdd_4_lut_25949 (.A(n30754), .B(n32470), .C(n1318), .D(n1286[3]), 
         .Z(n33741)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam n30754_bdd_4_lut_25949.init = 16'hee0f;
    FD1P3IX buffer_0___i22 (.D(n28240), .SP(n7986), .CD(n32395), .CK(debug_c_c), 
            .Q(\buffer[2] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i22.GSR = "ENABLED";
    LUT4 n30754_bdd_4_lut (.A(bufcount[1]), .B(n1286[4]), .C(bufcount[0]), 
         .D(bufcount[3]), .Z(n33743)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam n30754_bdd_4_lut.init = 16'h0080;
    FD1P3IX buffer_0___i23 (.D(n28251), .SP(n7986), .CD(n32395), .CK(debug_c_c), 
            .Q(\buffer[2] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i23.GSR = "ENABLED";
    FD1P3IX buffer_0___i24 (.D(n28228), .SP(n7986), .CD(n32395), .CK(debug_c_c), 
            .Q(\buffer[2] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i24.GSR = "ENABLED";
    FD1P3IX buffer_0___i25 (.D(n28323), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[3] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i25.GSR = "ENABLED";
    FD1P3IX buffer_0___i26 (.D(n28306), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[3] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i26.GSR = "ENABLED";
    FD1P3IX buffer_0___i27 (.D(n28197), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[3] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i27.GSR = "ENABLED";
    FD1P3IX buffer_0___i28 (.D(n28223), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[3] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i28.GSR = "ENABLED";
    FD1P3IX buffer_0___i29 (.D(n28297), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[3] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i29.GSR = "ENABLED";
    FD1P3IX buffer_0___i30 (.D(n28200), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[3] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i30.GSR = "ENABLED";
    FD1P3IX buffer_0___i31 (.D(n28206), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[3] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i31.GSR = "ENABLED";
    FD1P3IX buffer_0___i32 (.D(n28201), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[3] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i32.GSR = "ENABLED";
    FD1P3IX buffer_0___i33 (.D(n28204), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[4] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i33.GSR = "ENABLED";
    FD1P3IX buffer_0___i34 (.D(n28190), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[4] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i34.GSR = "ENABLED";
    FD1P3IX buffer_0___i35 (.D(n28344), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[4] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i35.GSR = "ENABLED";
    FD1P3IX buffer_0___i36 (.D(n28336), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[4] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i36.GSR = "ENABLED";
    FD1P3IX buffer_0___i37 (.D(n28343), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[4] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i37.GSR = "ENABLED";
    FD1P3IX buffer_0___i38 (.D(n28341), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[4] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i38.GSR = "ENABLED";
    FD1P3IX buffer_0___i39 (.D(n28338), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[4] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i39.GSR = "ENABLED";
    FD1P3IX buffer_0___i40 (.D(n28305), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[4] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i40.GSR = "ENABLED";
    FD1P3IX buffer_0___i41 (.D(n28358), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[5] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i41.GSR = "ENABLED";
    FD1P3IX buffer_0___i42 (.D(n28370), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[5] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i42.GSR = "ENABLED";
    FD1P3IX buffer_0___i43 (.D(n28184), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[5] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i43.GSR = "ENABLED";
    FD1P3IX buffer_0___i44 (.D(n28314), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[5] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i44.GSR = "ENABLED";
    FD1P3IX buffer_0___i45 (.D(n28283), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[5] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i45.GSR = "ENABLED";
    FD1P3IX buffer_0___i46 (.D(n28339), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[5] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i46.GSR = "ENABLED";
    FD1P3IX buffer_0___i47 (.D(n28303), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[5] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i47.GSR = "ENABLED";
    FD1P3IX buffer_0___i48 (.D(n28302), .SP(n7986), .CD(n34319), .CK(debug_c_c), 
            .Q(\buffer[5] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=57, LSE_LLINE=475, LSE_RLINE=485 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam buffer_0___i48.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_136 (.A(databus[26]), .B(n5_adj_72), .C(n1286[13]), 
         .D(n30202), .Z(n28184)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_136.init = 16'hffec;
    FD1P3AX rw_498_rep_422 (.D(n1286[10]), .SP(n2539), .CK(debug_c_c), 
            .Q(n34317));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam rw_498_rep_422.GSR = "ENABLED";
    LUT4 i461_2_lut (.A(n9), .B(n1304), .Z(n1398)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i461_2_lut.init = 16'h4444;
    LUT4 i7972_4_lut (.A(escape), .B(n11477), .C(n6_adj_73), .D(n1286[3]), 
         .Z(n9337)) /* synthesis lut_function=(!(A (C (D))+!A (B+!(C (D))))) */ ;
    defparam i7972_4_lut.init = 16'h1aaa;
    LUT4 i2_2_lut_adj_137 (.A(debug_c_7), .B(n32444), .Z(n6_adj_73)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_adj_137.init = 16'h8888;
    LUT4 select_1742_Select_42_i5_4_lut (.A(\buffer[5] [2]), .B(n1286[4]), 
         .C(rx_data[2]), .D(n30488), .Z(n5_adj_72)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_42_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_138 (.A(databus[27]), .B(n5_adj_74), .C(n1286[13]), 
         .D(n30203), .Z(n28314)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_138.init = 16'hffec;
    LUT4 select_1742_Select_43_i5_4_lut (.A(\buffer[5] [3]), .B(n1286[4]), 
         .C(rx_data[3]), .D(n30488), .Z(n5_adj_74)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_43_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_139 (.A(databus[28]), .B(n5_adj_75), .C(n1286[13]), 
         .D(n30204), .Z(n28283)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_139.init = 16'hffec;
    LUT4 i1_2_lut_adj_140 (.A(register_addr[1]), .B(\steps_reg[5]_adj_34 ), 
         .Z(n14_adj_35)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_140.init = 16'h8888;
    LUT4 select_1742_Select_44_i5_4_lut (.A(\buffer[5] [4]), .B(n1286[4]), 
         .C(rx_data[4]), .D(n30488), .Z(n5_adj_75)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_44_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_adj_141 (.A(register_addr[1]), .B(\steps_reg[3]_adj_36 ), 
         .Z(n15_adj_37)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_141.init = 16'h8888;
    PFUMX i25224 (.BLUT(n32271), .ALUT(n32266), .C0(n9), .Z(n32272));
    LUT4 i2_4_lut_adj_142 (.A(databus[0]), .B(n5_adj_80), .C(n1286[13]), 
         .D(n30183), .Z(n28255)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_142.init = 16'hffec;
    LUT4 i2_4_lut_adj_143 (.A(databus[29]), .B(n5_adj_81), .C(n1286[13]), 
         .D(n30206), .Z(n28339)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_143.init = 16'hffec;
    LUT4 i1_2_lut_adj_144 (.A(register_addr[1]), .B(\steps_reg[5]_adj_38 ), 
         .Z(n14_adj_39)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_144.init = 16'h8888;
    LUT4 select_1742_Select_16_i5_4_lut (.A(\buffer[2] [0]), .B(n1286[4]), 
         .C(rx_data[0]), .D(n30512), .Z(n5_adj_80)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_16_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_adj_145 (.A(register_addr[1]), .B(\steps_reg[3]_adj_40 ), 
         .Z(n15_adj_41)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_145.init = 16'h8888;
    LUT4 select_1742_Select_45_i5_4_lut (.A(\buffer[5] [5]), .B(n1286[4]), 
         .C(rx_data[5]), .D(n30488), .Z(n5_adj_81)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_45_i5_4_lut.init = 16'h88c0;
    LUT4 i1_2_lut_rep_419 (.A(n1286[6]), .B(n1286[11]), .Z(n32513)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_rep_419.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_146 (.A(n1286[6]), .B(n1286[11]), .C(n32444), 
         .Z(n18427)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_3_lut_adj_146.init = 16'he0e0;
    LUT4 i2_4_lut_adj_147 (.A(databus[30]), .B(n5_adj_86), .C(n1286[13]), 
         .D(n30199), .Z(n28303)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_147.init = 16'hffec;
    LUT4 mux_1314_i29_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[28]), 
         .D(n224[28]), .Z(n3181[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i29_3_lut_4_lut.init = 16'hf780;
    LUT4 i2882_2_lut_rep_421 (.A(\sendcount[1] ), .B(sendcount[0]), .Z(n32515)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i2882_2_lut_rep_421.init = 16'h9999;
    LUT4 n11281_bdd_4_lut_4_lut (.A(\sendcount[1] ), .B(sendcount[0]), .C(\buffer[5] [0]), 
         .D(\buffer[4] [0]), .Z(n32270)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam n11281_bdd_4_lut_4_lut.init = 16'h6420;
    LUT4 i13874_2_lut_2_lut_3_lut (.A(\sendcount[1] ), .B(sendcount[0]), 
         .C(n9_c), .Z(n19[1])) /* synthesis lut_function=(!(A (B (C))+!A !(B+!(C)))) */ ;
    defparam i13874_2_lut_2_lut_3_lut.init = 16'h6f6f;
    LUT4 i1_2_lut_3_lut_adj_148 (.A(rx_data[1]), .B(rx_data[4]), .C(rx_data[3]), 
         .Z(n11539)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(133[11] 166[18])
    defparam i1_2_lut_3_lut_adj_148.init = 16'h0808;
    LUT4 select_1742_Select_46_i5_4_lut (.A(\buffer[5] [6]), .B(n1286[4]), 
         .C(rx_data[6]), .D(n30488), .Z(n5_adj_86)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_46_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_149 (.A(n32380), .B(sendcount[3]), .C(n9_c), .D(n8679), 
         .Z(n28153)) /* synthesis lut_function=(!(A+(B ((D)+!C)+!B !(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i2_4_lut_adj_149.init = 16'h1040;
    LUT4 i2_4_lut_adj_150 (.A(databus[31]), .B(n5_adj_88), .C(n1286[13]), 
         .D(n30205), .Z(n28302)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_150.init = 16'hffec;
    LUT4 select_1742_Select_47_i5_4_lut (.A(\buffer[5] [7]), .B(n1286[4]), 
         .C(rx_data[7]), .D(n30488), .Z(n5_adj_88)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_47_i5_4_lut.init = 16'h88c0;
    LUT4 mux_1384_i1_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[0]), 
         .D(n224_adj_42[0]), .Z(n3451[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i1_3_lut_4_lut.init = 16'hf780;
    PFUMX i8317 (.BLUT(n14082), .ALUT(n1682[1]), .C0(n1687), .Z(n14083));
    PFUMX i7658 (.BLUT(n13423), .ALUT(n28389), .C0(n1687), .Z(n13424));
    LUT4 reduce_or_453_i1_3_lut_4_lut (.A(n32463), .B(n11639), .C(\buffer[0] [7]), 
         .D(n1286[9]), .Z(n1391)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(158[15] 160[18])
    defparam reduce_or_453_i1_3_lut_4_lut.init = 16'hff80;
    LUT4 mux_1384_i16_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[15]), 
         .D(n224_adj_42[15]), .Z(n3451[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1314_i1_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[0]), 
         .D(n224[0]), .Z(n3181[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_151 (.A(n1286[4]), .B(\buffer[0] [0]), .C(n11_adj_16), 
         .D(n14_adj_43), .Z(n29188)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_151.init = 16'heca0;
    LUT4 i2_3_lut (.A(n1286[19]), .B(n1286[16]), .C(n11238), .Z(n28369)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i2_3_lut.init = 16'hefef;
    LUT4 i24656_2_lut (.A(sendcount[0]), .B(n9_c), .Z(n20282)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i24656_2_lut.init = 16'h7777;
    LUT4 i1_4_lut_adj_152 (.A(sendcount[4]), .B(n1), .C(n6_adj_91), .D(n11271), 
         .Z(n9_c)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i1_4_lut_adj_152.init = 16'hfeff;
    LUT4 i24777_3_lut (.A(n32444), .B(n1286[20]), .C(n1286[17]), .Z(n11238)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i24777_3_lut.init = 16'h0202;
    LUT4 mux_1384_i15_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[14]), 
         .D(n224_adj_42[14]), .Z(n3451[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 equal_48_i1_3_lut (.A(sendcount[0]), .B(n5), .C(n6), .Z(n1)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam equal_48_i1_3_lut.init = 16'h5656;
    LUT4 i2_4_lut_adj_153 (.A(\reg_size[2] ), .B(sendcount[3]), .C(sendcount[2]), 
         .D(n32486), .Z(n6_adj_91)) /* synthesis lut_function=(A (B (C+!(D))+!B ((D)+!C))+!A (B+!(C (D)+!C !(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(268[12:39])
    defparam i2_4_lut_adj_153.init = 16'he7de;
    LUT4 mux_1578_i5_3_lut (.A(n9241[4]), .B(sendcount[0]), .C(n9), .Z(n4846[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1578_i5_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_4_i4_3_lut (.A(\buffer[4] [4]), .B(\buffer[5] [4]), 
         .C(sendcount[0]), .Z(n4_adj_26)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_4_i4_3_lut.init = 16'hacac;
    LUT4 mux_1578_i3_3_lut (.A(n9241[2]), .B(sendcount[0]), .C(n9), .Z(n4846[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1578_i3_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_2_i4_3_lut (.A(\buffer[4] [2]), .B(\buffer[5] [2]), 
         .C(sendcount[0]), .Z(n4_adj_25)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_2_i4_3_lut.init = 16'hacac;
    LUT4 i1_4_lut_adj_154 (.A(n1286[4]), .B(\buffer[1] [7]), .C(n11_adj_17), 
         .D(n14_adj_43), .Z(n29192)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_154.init = 16'heca0;
    LUT4 mux_1578_i2_3_lut (.A(n9241[1]), .B(sendcount[0]), .C(n9), .Z(n4846[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(249[9] 267[16])
    defparam mux_1578_i2_3_lut.init = 16'hcaca;
    LUT4 mux_429_Mux_1_i4_3_lut (.A(\buffer[4] [1]), .B(\buffer[5] [1]), 
         .C(sendcount[0]), .Z(n4_c)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(264[31:44])
    defparam mux_429_Mux_1_i4_3_lut.init = 16'hacac;
    LUT4 i5_4_lut_adj_155 (.A(n9_adj_53), .B(n1286[15]), .C(n8_adj_57), 
         .D(n1286[1]), .Z(debug_c_2)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i5_4_lut_adj_155.init = 16'hfffe;
    LUT4 i1_4_lut_adj_156 (.A(n1286[2]), .B(n32478), .C(n8_adj_95), .D(n1286[18]), 
         .Z(debug_c_3)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_156.init = 16'hfffe;
    LUT4 i3_4_lut_adj_157 (.A(n32482), .B(n1286[10]), .C(n4_adj_96), .D(n1286[6]), 
         .Z(n8_adj_95)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_157.init = 16'hfffe;
    LUT4 i1_2_lut_adj_158 (.A(n1286[11]), .B(n1286[7]), .Z(n4_adj_96)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_158.init = 16'heeee;
    LUT4 i4_4_lut_adj_159 (.A(n1286[20]), .B(n30537), .C(n32484), .D(n6_adj_97), 
         .Z(debug_c_4)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i4_4_lut_adj_159.init = 16'hfffe;
    LUT4 i1_2_lut_adj_160 (.A(n1286[4]), .B(n1286[6]), .Z(n6_adj_97)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam i1_2_lut_adj_160.init = 16'heeee;
    LUT4 i4_4_lut_adj_161 (.A(n1310), .B(n30537), .C(n32483), .D(n6_adj_98), 
         .Z(debug_c_5)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4_4_lut_adj_161.init = 16'hfffe;
    LUT4 i1_2_lut_adj_162 (.A(n1286[13]), .B(n1286[10]), .Z(n6_adj_98)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_2_lut_adj_162.init = 16'heeee;
    LUT4 mux_1314_i32_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[31]), 
         .D(n224[31]), .Z(n3181[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i32_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_163 (.A(n30390), .B(debug_c_7), .C(n1318), .D(n1286[1]), 
         .Z(n11936)) /* synthesis lut_function=(A+!(B+!(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_163.init = 16'hbbba;
    LUT4 i3_4_lut_adj_164 (.A(sendcount[3]), .B(n32476), .C(sendcount[2]), 
         .D(n32475), .Z(n30390)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_164.init = 16'h0200;
    LUT4 i2_4_lut_adj_165 (.A(databus[4]), .B(n5_adj_100), .C(n1286[13]), 
         .D(n30175), .Z(n28243)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_165.init = 16'hffec;
    LUT4 select_1742_Select_20_i5_4_lut (.A(\buffer[2] [4]), .B(n1286[4]), 
         .C(rx_data[4]), .D(n30512), .Z(n5_adj_100)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_20_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_166 (.A(databus[5]), .B(n5_adj_101), .C(n1286[13]), 
         .D(n30182), .Z(n28240)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_166.init = 16'hffec;
    LUT4 select_1742_Select_21_i5_4_lut (.A(\buffer[2] [5]), .B(n1286[4]), 
         .C(rx_data[5]), .D(n30512), .Z(n5_adj_101)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_21_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_167 (.A(databus[6]), .B(n5_adj_102), .C(n1286[13]), 
         .D(n30185), .Z(n28251)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_167.init = 16'hffec;
    LUT4 select_1742_Select_22_i5_4_lut (.A(\buffer[2] [6]), .B(n1286[4]), 
         .C(rx_data[6]), .D(n30512), .Z(n5_adj_102)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_22_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_168 (.A(databus[7]), .B(n5_adj_103), .C(n1286[13]), 
         .D(n30186), .Z(n28228)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_168.init = 16'hffec;
    LUT4 select_1742_Select_23_i5_4_lut (.A(\buffer[2] [7]), .B(n1286[4]), 
         .C(rx_data[7]), .D(n30512), .Z(n5_adj_103)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_23_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_169 (.A(databus[8]), .B(n5_adj_104), .C(n1286[13]), 
         .D(n30187), .Z(n28323)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_169.init = 16'hffec;
    LUT4 select_1742_Select_24_i5_4_lut (.A(\buffer[3] [0]), .B(n1286[4]), 
         .C(rx_data[0]), .D(n30511), .Z(n5_adj_104)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_24_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_170 (.A(databus[9]), .B(n5_adj_105), .C(n1286[13]), 
         .D(n30188), .Z(n28306)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_170.init = 16'hffec;
    LUT4 select_1742_Select_25_i5_4_lut (.A(\buffer[3] [1]), .B(n1286[4]), 
         .C(rx_data[1]), .D(n30511), .Z(n5_adj_105)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_25_i5_4_lut.init = 16'h88c0;
    LUT4 i24731_2_lut_2_lut (.A(n32444), .B(n7986), .Z(n12022)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i24731_2_lut_2_lut.init = 16'hdddd;
    LUT4 i2_4_lut_adj_171 (.A(databus[10]), .B(n5_adj_106), .C(n1286[13]), 
         .D(n30189), .Z(n28197)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_171.init = 16'hffec;
    LUT4 select_1742_Select_26_i5_4_lut (.A(\buffer[3] [2]), .B(n1286[4]), 
         .C(rx_data[2]), .D(n30511), .Z(n5_adj_106)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_26_i5_4_lut.init = 16'h88c0;
    LUT4 mux_1384_i14_3_lut_4_lut (.A(n30310), .B(n32343), .C(databus[13]), 
         .D(n224_adj_42[13]), .Z(n3451[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1384_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i24395_4_lut (.A(n30619), .B(rx_data[2]), .C(rx_data[1]), .D(n30734), 
         .Z(n30754)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24395_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_172 (.A(databus[11]), .B(n5_adj_108), .C(n1286[13]), 
         .D(n30193), .Z(n28223)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_172.init = 16'hffec;
    LUT4 i3_4_lut_adj_173 (.A(n34320), .B(n32503), .C(register_addr[2]), 
         .D(n30401), .Z(n11753)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i3_4_lut_adj_173.init = 16'h0100;
    LUT4 select_1742_Select_27_i5_4_lut (.A(\buffer[3] [3]), .B(n1286[4]), 
         .C(rx_data[3]), .D(n30511), .Z(n5_adj_108)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_27_i5_4_lut.init = 16'h88c0;
    LUT4 i24375_4_lut (.A(rx_data[4]), .B(rx_data[3]), .C(rx_data[0]), 
         .D(rx_data[1]), .Z(n30734)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i24375_4_lut.init = 16'hffef;
    LUT4 i24264_3_lut (.A(rx_data[6]), .B(rx_data[7]), .C(rx_data[5]), 
         .Z(n30619)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i24264_3_lut.init = 16'hfefe;
    LUT4 i24767_4_lut (.A(n7), .B(n30708), .C(n32470), .D(n1286[3]), 
         .Z(n7986)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C+!(D))))) */ ;
    defparam i24767_4_lut.init = 16'h0544;
    LUT4 i24349_3_lut (.A(n1286[13]), .B(n1318), .C(n1286[4]), .Z(n30708)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i24349_3_lut.init = 16'hfefe;
    LUT4 i2_4_lut_adj_174 (.A(databus[12]), .B(n5_adj_109), .C(n1286[13]), 
         .D(n30178), .Z(n28297)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_174.init = 16'hffec;
    LUT4 i4913_3_lut (.A(busy), .B(n1286[20]), .C(n1286[19]), .Z(n10677)) /* synthesis lut_function=(A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i4913_3_lut.init = 16'ha8a8;
    LUT4 select_1742_Select_28_i5_4_lut (.A(\buffer[3] [4]), .B(n1286[4]), 
         .C(rx_data[4]), .D(n30511), .Z(n5_adj_109)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_28_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_175 (.A(databus[13]), .B(n5_adj_110), .C(n1286[13]), 
         .D(n30192), .Z(n28200)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_175.init = 16'hffec;
    LUT4 select_1742_Select_29_i5_4_lut (.A(\buffer[3] [5]), .B(n1286[4]), 
         .C(rx_data[5]), .D(n30511), .Z(n5_adj_110)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_29_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut_adj_176 (.A(n1286[4]), .B(\buffer[1] [6]), .C(n11_adj_18), 
         .D(n14_adj_43), .Z(n29190)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_176.init = 16'heca0;
    LUT4 i2_4_lut_adj_177 (.A(databus[14]), .B(n5_adj_111), .C(n1286[13]), 
         .D(n30194), .Z(n28206)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_177.init = 16'hffec;
    LUT4 select_1742_Select_30_i5_4_lut (.A(\buffer[3] [6]), .B(n1286[4]), 
         .C(rx_data[6]), .D(n30511), .Z(n5_adj_111)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_30_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_178 (.A(databus[15]), .B(n5_adj_112), .C(n1286[13]), 
         .D(n30191), .Z(n28201)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_178.init = 16'hffec;
    LUT4 i1_4_lut_adj_179 (.A(n1286[4]), .B(\buffer[1] [5]), .C(n11_adj_19), 
         .D(n14_adj_43), .Z(n29174)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_179.init = 16'heca0;
    LUT4 mux_1314_i31_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[30]), 
         .D(n224[30]), .Z(n3181[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i31_3_lut_4_lut.init = 16'hf780;
    LUT4 select_1742_Select_31_i5_4_lut (.A(\buffer[3] [7]), .B(n1286[4]), 
         .C(rx_data[7]), .D(n30511), .Z(n5_adj_112)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_31_i5_4_lut.init = 16'h88c0;
    LUT4 i1_4_lut_adj_180 (.A(n1286[4]), .B(\buffer[1] [4]), .C(n11_adj_20), 
         .D(n14_adj_43), .Z(n29154)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_180.init = 16'heca0;
    LUT4 i1_4_lut_adj_181 (.A(n1286[4]), .B(\buffer[1] [3]), .C(n11_adj_21), 
         .D(n14_adj_43), .Z(n29264)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_181.init = 16'heca0;
    LUT4 i2_4_lut_adj_182 (.A(databus[3]), .B(n5_adj_114), .C(n1286[13]), 
         .D(n30179), .Z(n28238)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_182.init = 16'hffec;
    LUT4 i1_4_lut_adj_183 (.A(n1286[4]), .B(\buffer[1] [2]), .C(n11_adj_22), 
         .D(n14_adj_43), .Z(n29150)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_183.init = 16'heca0;
    LUT4 i14768_3_lut_rep_313 (.A(n1286[13]), .B(n32444), .C(n1304), .Z(n32407)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i14768_3_lut_rep_313.init = 16'hc8c8;
    LUT4 i2_4_lut_adj_184 (.A(databus[16]), .B(n5_adj_115), .C(n1286[13]), 
         .D(n30190), .Z(n28204)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_184.init = 16'hffec;
    LUT4 i3676_3_lut (.A(n1286[19]), .B(n1286[18]), .C(busy), .Z(n9437)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3676_3_lut.init = 16'hcece;
    LUT4 select_1742_Select_32_i5_4_lut (.A(\buffer[4] [0]), .B(n1286[4]), 
         .C(rx_data[0]), .D(n30487), .Z(n5_adj_115)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_32_i5_4_lut.init = 16'h88c0;
    LUT4 i24774_2_lut_3_lut_4_lut (.A(n1286[13]), .B(n32444), .C(n1304), 
         .D(n31948), .Z(n17)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;
    defparam i24774_2_lut_3_lut_4_lut.init = 16'hf700;
    LUT4 select_1742_Select_19_i5_4_lut (.A(\buffer[2] [3]), .B(n1286[4]), 
         .C(rx_data[3]), .D(n30512), .Z(n5_adj_114)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_19_i5_4_lut.init = 16'h88c0;
    LUT4 i24660_2_lut_rep_286_3_lut (.A(n1286[13]), .B(n32444), .C(n1304), 
         .Z(n32380)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i24660_2_lut_rep_286_3_lut.init = 16'h0808;
    LUT4 i2_4_lut_adj_185 (.A(databus[17]), .B(n5_adj_116), .C(n1286[13]), 
         .D(n30181), .Z(n28190)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_185.init = 16'hffec;
    LUT4 select_1742_Select_33_i5_4_lut (.A(\buffer[4] [1]), .B(n1286[4]), 
         .C(rx_data[1]), .D(n30487), .Z(n5_adj_116)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_33_i5_4_lut.init = 16'h88c0;
    LUT4 i2_4_lut_adj_186 (.A(n38), .B(busy), .C(n31399), .D(n1286[17]), 
         .Z(n29350)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_186.init = 16'hfbfa;
    LUT4 i1_4_lut_adj_187 (.A(n1286[4]), .B(\buffer[1] [1]), .C(n11_adj_23), 
         .D(n14_adj_43), .Z(n29196)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_187.init = 16'heca0;
    LUT4 i1_4_lut_adj_188 (.A(n1286[15]), .B(esc_data[7]), .C(n8_adj_117), 
         .D(esc_data[0]), .Z(n38)) /* synthesis lut_function=(A (B+(C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_188.init = 16'ha8aa;
    LUT4 i3_4_lut_adj_189 (.A(n35), .B(esc_data[5]), .C(n55), .D(esc_data[6]), 
         .Z(n8_adj_117)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i3_4_lut_adj_189.init = 16'hfffe;
    LUT4 i2_4_lut_adj_190 (.A(databus[18]), .B(n5_adj_118), .C(n1286[13]), 
         .D(n30195), .Z(n28344)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_190.init = 16'hffec;
    LUT4 rx_data_2__bdd_4_lut (.A(rx_data[2]), .B(rx_data[3]), .C(rx_data[4]), 
         .D(rx_data[1]), .Z(n31474)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D))+!B !(C+(D))))) */ ;
    defparam rx_data_2__bdd_4_lut.init = 16'h6001;
    LUT4 i1_4_lut_adj_191 (.A(n1286[4]), .B(\buffer[1] [0]), .C(n11_adj_24), 
         .D(n14_adj_43), .Z(n29200)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_191.init = 16'heca0;
    LUT4 select_1742_Select_34_i5_4_lut (.A(\buffer[4] [2]), .B(n1286[4]), 
         .C(rx_data[2]), .D(n30487), .Z(n5_adj_118)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_34_i5_4_lut.init = 16'h88c0;
    PFUMX i25279 (.BLUT(n32546), .ALUT(n32547), .C0(n32445), .Z(n32548));
    PFUMX i25277 (.BLUT(n32543), .ALUT(n32544), .C0(sendcount[0]), .Z(n32545));
    LUT4 i1_4_lut_adj_192 (.A(n1286[4]), .B(\buffer[0] [7]), .C(n11), 
         .D(n14_adj_43), .Z(n29152)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i1_4_lut_adj_192.init = 16'heca0;
    PFUMX i25275 (.BLUT(n32540), .ALUT(n32541), .C0(sendcount[0]), .Z(n32542));
    LUT4 i2_4_lut_adj_193 (.A(databus[2]), .B(n5_adj_119), .C(n1286[13]), 
         .D(n30184), .Z(n28252)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam i2_4_lut_adj_193.init = 16'hffec;
    PFUMX i25273 (.BLUT(n32537), .ALUT(n32538), .C0(sendcount[0]), .Z(n32539));
    LUT4 mux_1314_i30_3_lut_4_lut (.A(n32358), .B(n30258), .C(databus[29]), 
         .D(n224[29]), .Z(n3181[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(72[9] 328[6])
    defparam mux_1314_i30_3_lut_4_lut.init = 16'hf780;
    PFUMX i25271 (.BLUT(n32534), .ALUT(n32535), .C0(sendcount[0]), .Z(n32536));
    PFUMX i25269 (.BLUT(n32531), .ALUT(n32532), .C0(sendcount[0]), .Z(n32533));
    PFUMX i25267 (.BLUT(n32528), .ALUT(n32529), .C0(sendcount[0]), .Z(n32530));
    PFUMX i25265 (.BLUT(n32525), .ALUT(n32526), .C0(sendcount[0]), .Z(n32527));
    PFUMX i25263 (.BLUT(n32522), .ALUT(n32523), .C0(sendcount[0]), .Z(n32524));
    LUT4 select_1742_Select_18_i5_4_lut (.A(\buffer[2] [2]), .B(n1286[4]), 
         .C(rx_data[2]), .D(n30512), .Z(n5_adj_119)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(89[6] 326[13])
    defparam select_1742_Select_18_i5_4_lut.init = 16'h88c0;
    \UARTTransmitter(baud_div=12)  uart_output (.\reset_count[14] (\reset_count[14] ), 
            .\reset_count[12] (\reset_count[12] ), .\reset_count[13] (\reset_count[13] ), 
            .n32444(n32444), .n32395(n32395), .tx_data({tx_data}), .send(send), 
            .\reset_count[11] (\reset_count[11] ), .n19877(n19877), .\reset_count[8] (\reset_count[8] ), 
            .n27962(n27962), .busy(busy), .n34319(n34319), .n9395(n9395), 
            .\reset_count[10] (\reset_count[10] ), .\reset_count[9] (\reset_count[9] ), 
            .debug_c_c(debug_c_c), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(65[30] 70[52])
    \UARTReceiver(baud_div=12)  uart_input (.state({state}), .n32(n32), 
            .rdata({Open_46, Open_47, Open_48, Open_49, Open_50, Open_51, 
            Open_52, \rdata[0] }), .debug_c_c(debug_c_c), .n32444(n32444), 
            .bclk(bclk), .rx_data({rx_data}), .n32395(n32395), .n34319(n34319), 
            .n29158(n29158), .\rdata[1] (\rdata[1] ), .n9396_c(n9396_c), 
            .n31442(n31442), .debug_c_7(debug_c_7), .n183(n183), .n31427(n31427), 
            .n32432(n32432), .n32409(n32409), .n32495(n32495), .n32494(n32494), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(60[27] 64[39])
    
endmodule
//
// Verilog Description of module \UARTTransmitter(baud_div=12) 
//

module \UARTTransmitter(baud_div=12)  (\reset_count[14] , \reset_count[12] , 
            \reset_count[13] , n32444, n32395, tx_data, send, \reset_count[11] , 
            n19877, \reset_count[8] , n27962, busy, n34319, n9395, 
            \reset_count[10] , \reset_count[9] , debug_c_c, GND_net) /* synthesis syn_module_defined=1 */ ;
    input \reset_count[14] ;
    input \reset_count[12] ;
    input \reset_count[13] ;
    output n32444;
    output n32395;
    input [7:0]tx_data;
    input send;
    input \reset_count[11] ;
    output n19877;
    input \reset_count[8] ;
    input n27962;
    output busy;
    output n34319;
    output n9395;
    input \reset_count[10] ;
    input \reset_count[9] ;
    input debug_c_c;
    input GND_net;
    
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n30400, n7, n10;
    wire [3:0]state;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(102[12:17])
    
    wire n104, n31425;
    wire [7:0]tdata;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(101[12:17])
    
    wire n7984, n12208, n29048, n17, n17_adj_9, n31424, n30827, 
        n30828, n30829, n31936, n13675, n31423, n31935, n30386, 
        n30385, n32400, n2533, n30231, n19754, n2;
    
    LUT4 i1_4_lut_rep_350 (.A(\reset_count[14] ), .B(\reset_count[12] ), 
         .C(\reset_count[13] ), .D(n30400), .Z(n32444)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_rep_350.init = 16'hfaea;
    LUT4 i14745_1_lut_rep_301_4_lut (.A(\reset_count[14] ), .B(\reset_count[12] ), 
         .C(\reset_count[13] ), .D(n30400), .Z(n32395)) /* synthesis lut_function=(!(A+(B (C)+!B (C (D))))) */ ;
    defparam i14745_1_lut_rep_301_4_lut.init = 16'h0515;
    PFUMX Mux_22_i15 (.BLUT(n7), .ALUT(n10), .C0(state[3]), .Z(n104)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;
    FD1S3IX state__i0 (.D(n31425), .CK(bclk), .CD(n32395), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i0.GSR = "ENABLED";
    FD1P3AX tdata_i0_i0 (.D(tx_data[0]), .SP(n7984), .CK(bclk), .Q(tdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i0.GSR = "ENABLED";
    FD1P3AX tdata_i0_i7 (.D(tx_data[7]), .SP(n7984), .CK(bclk), .Q(tdata[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i7.GSR = "ENABLED";
    FD1P3AX tdata_i0_i6 (.D(tx_data[6]), .SP(n7984), .CK(bclk), .Q(tdata[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i6.GSR = "ENABLED";
    FD1P3AX tdata_i0_i5 (.D(tx_data[5]), .SP(n7984), .CK(bclk), .Q(tdata[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i5.GSR = "ENABLED";
    FD1P3AX tdata_i0_i4 (.D(tx_data[4]), .SP(n7984), .CK(bclk), .Q(tdata[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i4.GSR = "ENABLED";
    FD1P3AX tdata_i0_i3 (.D(tx_data[3]), .SP(n7984), .CK(bclk), .Q(tdata[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i3.GSR = "ENABLED";
    FD1P3AX tdata_i0_i2 (.D(tx_data[2]), .SP(n7984), .CK(bclk), .Q(tdata[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i2.GSR = "ENABLED";
    FD1P3AX tdata_i0_i1 (.D(tx_data[1]), .SP(n7984), .CK(bclk), .Q(tdata[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tdata_i0_i1.GSR = "ENABLED";
    FD1P3AX state__i3 (.D(n29048), .SP(n12208), .CK(bclk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i3.GSR = "ENABLED";
    LUT4 i27_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), .D(state[3]), 
         .Z(n17)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B !(C+(D))))) */ ;
    defparam i27_4_lut_4_lut.init = 16'h15fe;
    LUT4 i24_4_lut_4_lut (.A(state[3]), .B(state[0]), .C(state[1]), .D(send), 
         .Z(n17_adj_9)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;
    defparam i24_4_lut_4_lut.init = 16'h8001;
    LUT4 i2_4_lut (.A(\reset_count[11] ), .B(n19877), .C(\reset_count[8] ), 
         .D(n27962), .Z(n30400)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 state_1__bdd_4_lut (.A(state[1]), .B(state[3]), .C(state[0]), 
         .D(send), .Z(n31424)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(B (C)+!B (C+!(D)))) */ ;
    defparam state_1__bdd_4_lut.init = 16'h8f0e;
    PFUMX i24470 (.BLUT(n30827), .ALUT(n30828), .C0(state[1]), .Z(n30829));
    FD1P3IX busy_34 (.D(n13675), .SP(n31936), .CD(n34319), .CK(bclk), 
            .Q(busy));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam busy_34.GSR = "ENABLED";
    LUT4 state_1__bdd_2_lut (.A(state[3]), .B(state[0]), .Z(n31423)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam state_1__bdd_2_lut.init = 16'h1111;
    LUT4 state_2__bdd_4_lut_25786 (.A(state[0]), .B(state[3]), .C(state[1]), 
         .D(send), .Z(n31935)) /* synthesis lut_function=(A (B (C))+!A !(B+(C+!(D)))) */ ;
    defparam state_2__bdd_4_lut_25786.init = 16'h8180;
    LUT4 n31935_bdd_2_lut (.A(n31935), .B(state[2]), .Z(n31936)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n31935_bdd_2_lut.init = 16'h2222;
    LUT4 i14745_1_lut_rep_424 (.A(\reset_count[14] ), .B(\reset_count[12] ), 
         .C(\reset_count[13] ), .D(n30400), .Z(n34319)) /* synthesis lut_function=(!(A+(B (C)+!B (C (D))))) */ ;
    defparam i14745_1_lut_rep_424.init = 16'h0515;
    FD1P3AX state__i1 (.D(n30386), .SP(n12208), .CK(bclk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i1.GSR = "ENABLED";
    FD1P3AX state__i2 (.D(n30385), .SP(n12208), .CK(bclk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam state__i2.GSR = "ENABLED";
    FD1P3JX tx_35 (.D(n104), .SP(n17), .PD(n32395), .CK(bclk), .Q(n9395)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=30, LSE_RCOL=52, LSE_LLINE=65, LSE_RLINE=70 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam tx_35.GSR = "ENABLED";
    LUT4 i24468_3_lut (.A(tdata[2]), .B(tdata[3]), .C(state[0]), .Z(n30827)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24468_3_lut.init = 16'hcaca;
    LUT4 i24469_3_lut (.A(tdata[4]), .B(tdata[5]), .C(state[0]), .Z(n30828)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24469_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(\reset_count[10] ), .B(\reset_count[9] ), .Z(n19877)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i3_1_lut (.A(state[3]), .Z(n13675)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i3_1_lut.init = 16'h5555;
    LUT4 i1_3_lut (.A(state[1]), .B(n32400), .C(state[0]), .Z(n30386)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4848;
    LUT4 i1_2_lut_adj_49 (.A(state[0]), .B(state[1]), .Z(n2533)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_49.init = 16'h8888;
    LUT4 i2_4_lut_adj_50 (.A(n30231), .B(state[2]), .C(n19754), .D(n32444), 
         .Z(n7984)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i2_4_lut_adj_50.init = 16'h0200;
    LUT4 i1_2_lut_adj_51 (.A(send), .B(state[3]), .Z(n30231)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_51.init = 16'h2222;
    LUT4 i14022_2_lut (.A(state[1]), .B(state[0]), .Z(n19754)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14022_2_lut.init = 16'heeee;
    LUT4 i24785_3_lut (.A(n32444), .B(n17_adj_9), .C(state[2]), .Z(n12208)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i24785_3_lut.init = 16'hf7f7;
    LUT4 i1_4_lut (.A(n32444), .B(state[3]), .C(state[2]), .D(n2533), 
         .Z(n29048)) /* synthesis lut_function=(!((B (C)+!B !(C (D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(107[9] 190[6])
    defparam i1_4_lut.init = 16'h2808;
    LUT4 i1_3_lut_rep_306 (.A(n32444), .B(state[2]), .C(state[3]), .Z(n32400)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i1_3_lut_rep_306.init = 16'h2a2a;
    LUT4 i1_3_lut_4_lut (.A(n32444), .B(state[2]), .C(state[3]), .D(n2533), 
         .Z(n30385)) /* synthesis lut_function=(!((B (C+(D))+!B !(D))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h2208;
    PFUMX i24900 (.BLUT(n31424), .ALUT(n31423), .C0(state[2]), .Z(n31425));
    LUT4 Mux_22_i7_4_lut (.A(n2), .B(n30829), .C(state[2]), .D(state[1]), 
         .Z(n7)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i7_4_lut.init = 16'hcac0;
    LUT4 Mux_22_i2_3_lut (.A(tdata[0]), .B(tdata[1]), .C(state[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i14259_4_lut (.A(tdata[6]), .B(state[1]), .C(tdata[7]), .D(state[0]), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(117[6] 188[13])
    defparam i14259_4_lut.init = 16'hfcee;
    \ClockDividerP(factor=12)  baud_gen (.debug_c_c(debug_c_c), .bclk(bclk), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(104[28] 106[50])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12) 
//

module \ClockDividerP(factor=12)  (debug_c_c, bclk, GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    output bclk;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    wire bclk /* synthesis SET_AS_NETWORK=\protocol_interface/uart_output/bclk */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(100[7:11])
    
    wire n55;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    
    wire n56, n4, n14394, n52, n44, n35, n54, n48, n36, n46, 
        n32, n50, n40;
    wire [31:0]n102;
    
    wire n7264, n27506, n27507, n27893, n27892, n27891, n27890, 
        n27889, n27888, n27887, n27886, n27885, n27884, n27883, 
        n27882, n27881, n27880, n27879, n27878, n27521, n27520, 
        n27519, n27518, n27517, n27516, n27515, n27514, n27513, 
        n27512, n27511, n27510, n27509, n27508;
    
    LUT4 i24755_4_lut (.A(n55), .B(count[1]), .C(n56), .D(n4), .Z(n14394)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i24755_4_lut.init = 16'h0400;
    LUT4 i26_4_lut (.A(count[14]), .B(n52), .C(n44), .D(count[6]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i27_4_lut (.A(n35), .B(n54), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(count[3]), .B(count[0]), .Z(n4)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i23_4_lut (.A(count[24]), .B(n46), .C(n32), .D(count[16]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i15_3_lut (.A(count[15]), .B(count[31]), .C(count[5]), .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i17_4_lut (.A(count[26]), .B(count[12]), .C(count[28]), .D(count[18]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[13]), .B(count[22]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(count[20]), .B(count[4]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i25_4_lut (.A(count[25]), .B(n50), .C(n40), .D(count[9]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(count[7]), .B(count[19]), .C(count[11]), .D(count[21]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[8]), .B(count[29]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i21_4_lut (.A(count[2]), .B(count[27]), .C(count[23]), .D(count[30]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i11_2_lut (.A(count[10]), .B(count[17]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam i11_2_lut.init = 16'heeee;
    FD1S3IX count_2181__i0 (.D(n102[0]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i0.GSR = "ENABLED";
    FD1S3AX clk_o_14 (.D(n7264), .CK(debug_c_c), .Q(bclk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=28, LSE_RCOL=50, LSE_LLINE=104, LSE_RLINE=106 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    CCU2D sub_1736_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27506), .COUT(n27507));
    defparam sub_1736_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_1736_add_2_4.INIT1 = 16'h5555;
    defparam sub_1736_add_2_4.INJECT1_0 = "NO";
    defparam sub_1736_add_2_4.INJECT1_1 = "NO";
    FD1S3IX count_2181__i1 (.D(n102[1]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i1.GSR = "ENABLED";
    FD1S3IX count_2181__i2 (.D(n102[2]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i2.GSR = "ENABLED";
    FD1S3IX count_2181__i3 (.D(n102[3]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i3.GSR = "ENABLED";
    FD1S3IX count_2181__i4 (.D(n102[4]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i4.GSR = "ENABLED";
    FD1S3IX count_2181__i5 (.D(n102[5]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i5.GSR = "ENABLED";
    FD1S3IX count_2181__i6 (.D(n102[6]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i6.GSR = "ENABLED";
    FD1S3IX count_2181__i7 (.D(n102[7]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i7.GSR = "ENABLED";
    FD1S3IX count_2181__i8 (.D(n102[8]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i8.GSR = "ENABLED";
    FD1S3IX count_2181__i9 (.D(n102[9]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i9.GSR = "ENABLED";
    FD1S3IX count_2181__i10 (.D(n102[10]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i10.GSR = "ENABLED";
    FD1S3IX count_2181__i11 (.D(n102[11]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i11.GSR = "ENABLED";
    FD1S3IX count_2181__i12 (.D(n102[12]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i12.GSR = "ENABLED";
    FD1S3IX count_2181__i13 (.D(n102[13]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i13.GSR = "ENABLED";
    FD1S3IX count_2181__i14 (.D(n102[14]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i14.GSR = "ENABLED";
    FD1S3IX count_2181__i15 (.D(n102[15]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i15.GSR = "ENABLED";
    FD1S3IX count_2181__i16 (.D(n102[16]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i16.GSR = "ENABLED";
    FD1S3IX count_2181__i17 (.D(n102[17]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i17.GSR = "ENABLED";
    FD1S3IX count_2181__i18 (.D(n102[18]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i18.GSR = "ENABLED";
    FD1S3IX count_2181__i19 (.D(n102[19]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i19.GSR = "ENABLED";
    FD1S3IX count_2181__i20 (.D(n102[20]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i20.GSR = "ENABLED";
    FD1S3IX count_2181__i21 (.D(n102[21]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i21.GSR = "ENABLED";
    FD1S3IX count_2181__i22 (.D(n102[22]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i22.GSR = "ENABLED";
    FD1S3IX count_2181__i23 (.D(n102[23]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i23.GSR = "ENABLED";
    FD1S3IX count_2181__i24 (.D(n102[24]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i24.GSR = "ENABLED";
    FD1S3IX count_2181__i25 (.D(n102[25]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i25.GSR = "ENABLED";
    FD1S3IX count_2181__i26 (.D(n102[26]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i26.GSR = "ENABLED";
    FD1S3IX count_2181__i27 (.D(n102[27]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i27.GSR = "ENABLED";
    FD1S3IX count_2181__i28 (.D(n102[28]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i28.GSR = "ENABLED";
    FD1S3IX count_2181__i29 (.D(n102[29]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i29.GSR = "ENABLED";
    FD1S3IX count_2181__i30 (.D(n102[30]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i30.GSR = "ENABLED";
    FD1S3IX count_2181__i31 (.D(n102[31]), .CK(debug_c_c), .CD(n14394), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181__i31.GSR = "ENABLED";
    CCU2D sub_1736_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27506));
    defparam sub_1736_add_2_2.INIT0 = 16'h0000;
    defparam sub_1736_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_1736_add_2_2.INJECT1_0 = "NO";
    defparam sub_1736_add_2_2.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27893), .S0(n102[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_33.INIT1 = 16'h0000;
    defparam count_2181_add_4_33.INJECT1_0 = "NO";
    defparam count_2181_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27892), .COUT(n27893), .S0(n102[29]), 
          .S1(n102[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_31.INJECT1_0 = "NO";
    defparam count_2181_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27891), .COUT(n27892), .S0(n102[27]), 
          .S1(n102[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_29.INJECT1_0 = "NO";
    defparam count_2181_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27890), .COUT(n27891), .S0(n102[25]), 
          .S1(n102[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_27.INJECT1_0 = "NO";
    defparam count_2181_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27889), .COUT(n27890), .S0(n102[23]), 
          .S1(n102[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_25.INJECT1_0 = "NO";
    defparam count_2181_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27888), .COUT(n27889), .S0(n102[21]), 
          .S1(n102[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_23.INJECT1_0 = "NO";
    defparam count_2181_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27887), .COUT(n27888), .S0(n102[19]), 
          .S1(n102[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_21.INJECT1_0 = "NO";
    defparam count_2181_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27886), .COUT(n27887), .S0(n102[17]), 
          .S1(n102[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_19.INJECT1_0 = "NO";
    defparam count_2181_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27885), .COUT(n27886), .S0(n102[15]), 
          .S1(n102[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_17.INJECT1_0 = "NO";
    defparam count_2181_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27884), .COUT(n27885), .S0(n102[13]), 
          .S1(n102[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_15.INJECT1_0 = "NO";
    defparam count_2181_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27883), .COUT(n27884), .S0(n102[11]), 
          .S1(n102[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_13.INJECT1_0 = "NO";
    defparam count_2181_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27882), .COUT(n27883), .S0(n102[9]), .S1(n102[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_11.INJECT1_0 = "NO";
    defparam count_2181_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27881), .COUT(n27882), .S0(n102[7]), .S1(n102[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_9.INJECT1_0 = "NO";
    defparam count_2181_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27880), .COUT(n27881), .S0(n102[5]), .S1(n102[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_7.INJECT1_0 = "NO";
    defparam count_2181_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27879), .COUT(n27880), .S0(n102[3]), .S1(n102[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_5.INJECT1_0 = "NO";
    defparam count_2181_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27878), .COUT(n27879), .S0(n102[1]), .S1(n102[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2181_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2181_add_4_3.INJECT1_0 = "NO";
    defparam count_2181_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2181_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27878), .S1(n102[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2181_add_4_1.INIT0 = 16'hF000;
    defparam count_2181_add_4_1.INIT1 = 16'h0555;
    defparam count_2181_add_4_1.INJECT1_0 = "NO";
    defparam count_2181_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27521), .S0(n7264));
    defparam sub_1736_add_2_cout.INIT0 = 16'h0000;
    defparam sub_1736_add_2_cout.INIT1 = 16'h0000;
    defparam sub_1736_add_2_cout.INJECT1_0 = "NO";
    defparam sub_1736_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27520), .COUT(n27521));
    defparam sub_1736_add_2_32.INIT0 = 16'h5555;
    defparam sub_1736_add_2_32.INIT1 = 16'h5555;
    defparam sub_1736_add_2_32.INJECT1_0 = "NO";
    defparam sub_1736_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27519), .COUT(n27520));
    defparam sub_1736_add_2_30.INIT0 = 16'h5555;
    defparam sub_1736_add_2_30.INIT1 = 16'h5555;
    defparam sub_1736_add_2_30.INJECT1_0 = "NO";
    defparam sub_1736_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27518), .COUT(n27519));
    defparam sub_1736_add_2_28.INIT0 = 16'h5555;
    defparam sub_1736_add_2_28.INIT1 = 16'h5555;
    defparam sub_1736_add_2_28.INJECT1_0 = "NO";
    defparam sub_1736_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27517), .COUT(n27518));
    defparam sub_1736_add_2_26.INIT0 = 16'h5555;
    defparam sub_1736_add_2_26.INIT1 = 16'h5555;
    defparam sub_1736_add_2_26.INJECT1_0 = "NO";
    defparam sub_1736_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27516), .COUT(n27517));
    defparam sub_1736_add_2_24.INIT0 = 16'h5555;
    defparam sub_1736_add_2_24.INIT1 = 16'h5555;
    defparam sub_1736_add_2_24.INJECT1_0 = "NO";
    defparam sub_1736_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27515), .COUT(n27516));
    defparam sub_1736_add_2_22.INIT0 = 16'h5555;
    defparam sub_1736_add_2_22.INIT1 = 16'h5555;
    defparam sub_1736_add_2_22.INJECT1_0 = "NO";
    defparam sub_1736_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27514), .COUT(n27515));
    defparam sub_1736_add_2_20.INIT0 = 16'h5555;
    defparam sub_1736_add_2_20.INIT1 = 16'h5555;
    defparam sub_1736_add_2_20.INJECT1_0 = "NO";
    defparam sub_1736_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27513), .COUT(n27514));
    defparam sub_1736_add_2_18.INIT0 = 16'h5555;
    defparam sub_1736_add_2_18.INIT1 = 16'h5555;
    defparam sub_1736_add_2_18.INJECT1_0 = "NO";
    defparam sub_1736_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27512), .COUT(n27513));
    defparam sub_1736_add_2_16.INIT0 = 16'h5555;
    defparam sub_1736_add_2_16.INIT1 = 16'h5555;
    defparam sub_1736_add_2_16.INJECT1_0 = "NO";
    defparam sub_1736_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27511), .COUT(n27512));
    defparam sub_1736_add_2_14.INIT0 = 16'h5555;
    defparam sub_1736_add_2_14.INIT1 = 16'h5555;
    defparam sub_1736_add_2_14.INJECT1_0 = "NO";
    defparam sub_1736_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27510), .COUT(n27511));
    defparam sub_1736_add_2_12.INIT0 = 16'h5555;
    defparam sub_1736_add_2_12.INIT1 = 16'h5555;
    defparam sub_1736_add_2_12.INJECT1_0 = "NO";
    defparam sub_1736_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27509), .COUT(n27510));
    defparam sub_1736_add_2_10.INIT0 = 16'h5555;
    defparam sub_1736_add_2_10.INIT1 = 16'h5555;
    defparam sub_1736_add_2_10.INJECT1_0 = "NO";
    defparam sub_1736_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27508), .COUT(n27509));
    defparam sub_1736_add_2_8.INIT0 = 16'h5555;
    defparam sub_1736_add_2_8.INIT1 = 16'h5555;
    defparam sub_1736_add_2_8.INJECT1_0 = "NO";
    defparam sub_1736_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_1736_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27507), .COUT(n27508));
    defparam sub_1736_add_2_6.INIT0 = 16'h5555;
    defparam sub_1736_add_2_6.INIT1 = 16'h5555;
    defparam sub_1736_add_2_6.INJECT1_0 = "NO";
    defparam sub_1736_add_2_6.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \UARTReceiver(baud_div=12) 
//

module \UARTReceiver(baud_div=12)  (state, n32, rdata, debug_c_c, n32444, 
            bclk, rx_data, n32395, n34319, n29158, \rdata[1] , n9396_c, 
            n31442, debug_c_7, n183, n31427, n32432, n32409, n32495, 
            n32494, GND_net) /* synthesis syn_module_defined=1 */ ;
    output [5:0]state;
    output n32;
    output [7:0]rdata;
    input debug_c_c;
    input n32444;
    output bclk;
    output [7:0]rx_data;
    input n32395;
    input n34319;
    input n29158;
    output \rdata[1] ;
    input n9396_c;
    input n31442;
    output debug_c_7;
    input n183;
    input n31427;
    input n32432;
    input n32409;
    input n32495;
    input n32494;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n29, n13984, n13985, n21, n17, n29092, n21_adj_7, n23, 
        n28810, n32449, n7934, n29228, n32493, n4, n7936, n31418;
    wire [5:0]n1;
    
    wire baud_reset, n29398, n31420, n7976, n7974, n7972, n7970, 
        n7968, n7966, n7964;
    wire [7:0]rdata_c;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(22[12:17])
    
    wire n7962, n7960, n7958, n7956, n7954, n7952, n7950, n32450, 
        n31419, n11696;
    wire [7:0]n78;
    
    wire n13, n11875, n30516, n29148, n4_adj_8, n19, n55, n27961, 
        n56, n2687, n23288, n219, n30483;
    
    PFUMX i8219 (.BLUT(n29), .ALUT(n13984), .C0(state[0]), .Z(n13985));
    PFUMX i32 (.BLUT(n21), .ALUT(n17), .C0(state[0]), .Z(n29092));
    PFUMX i36 (.BLUT(n21_adj_7), .ALUT(n23), .C0(state[5]), .Z(n28810));
    LUT4 i1_2_lut_rep_355 (.A(state[5]), .B(n32), .Z(n32449)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_2_lut_rep_355.init = 16'h4444;
    FD1P3AX rdata_i0_i0 (.D(n7934), .SP(n32444), .CK(debug_c_c), .Q(rdata[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i0.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut (.A(state[5]), .B(n32), .C(state[0]), .D(bclk), 
         .Z(n29228)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_3_lut_4_lut.init = 16'hf400;
    LUT4 i1_2_lut_3_lut (.A(state[3]), .B(n32493), .C(state[4]), .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    FD1P3AX data_i0_i0 (.D(n7936), .SP(n32444), .CK(debug_c_c), .Q(rx_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i0.GSR = "ENABLED";
    FD1S3IX state__i0 (.D(n29228), .CK(debug_c_c), .CD(n32395), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i0.GSR = "ENABLED";
    LUT4 n30396_bdd_3_lut_4_lut (.A(state[3]), .B(n32493), .C(bclk), .D(state[4]), 
         .Z(n31418)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;
    defparam n30396_bdd_3_lut_4_lut.init = 16'hf708;
    LUT4 mux_8_i4_3_lut_3_lut (.A(state[3]), .B(n32493), .C(bclk), .Z(n1[3])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;
    defparam mux_8_i4_3_lut_3_lut.init = 16'h6a6a;
    FD1S3JX baud_reset_52 (.D(n29398), .CK(debug_c_c), .PD(n32395), .Q(baud_reset)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam baud_reset_52.GSR = "ENABLED";
    LUT4 i8218_3_lut_3_lut (.A(state[3]), .B(n32493), .C(bclk), .Z(n13984)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;
    defparam i8218_3_lut_3_lut.init = 16'ha6a6;
    FD1S3IX state__i5 (.D(n28810), .CK(debug_c_c), .CD(n32395), .Q(state[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i5.GSR = "ENABLED";
    FD1S3IX state__i4 (.D(n31420), .CK(debug_c_c), .CD(n32395), .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i4.GSR = "ENABLED";
    FD1S3IX state__i3 (.D(n13985), .CK(debug_c_c), .CD(n34319), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i3.GSR = "ENABLED";
    FD1S3IX state__i2 (.D(n29092), .CK(debug_c_c), .CD(n34319), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i2.GSR = "ENABLED";
    FD1S3IX state__i1 (.D(n29158), .CK(debug_c_c), .CD(n34319), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam state__i1.GSR = "ENABLED";
    FD1P3AX data_i0_i7 (.D(n7976), .SP(n32444), .CK(debug_c_c), .Q(rx_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i7.GSR = "ENABLED";
    FD1P3AX data_i0_i6 (.D(n7974), .SP(n32444), .CK(debug_c_c), .Q(rx_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i6.GSR = "ENABLED";
    FD1P3AX data_i0_i5 (.D(n7972), .SP(n32444), .CK(debug_c_c), .Q(rx_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i5.GSR = "ENABLED";
    FD1P3AX data_i0_i4 (.D(n7970), .SP(n32444), .CK(debug_c_c), .Q(rx_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i4.GSR = "ENABLED";
    FD1P3AX data_i0_i3 (.D(n7968), .SP(n32444), .CK(debug_c_c), .Q(rx_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i3.GSR = "ENABLED";
    FD1P3AX data_i0_i2 (.D(n7966), .SP(n32444), .CK(debug_c_c), .Q(rx_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i2.GSR = "ENABLED";
    FD1P3AX data_i0_i1 (.D(n7964), .SP(n32444), .CK(debug_c_c), .Q(rx_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam data_i0_i1.GSR = "ENABLED";
    FD1P3AX rdata_i0_i7 (.D(n7962), .SP(n32444), .CK(debug_c_c), .Q(rdata_c[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i7.GSR = "ENABLED";
    FD1P3AX rdata_i0_i6 (.D(n7960), .SP(n32444), .CK(debug_c_c), .Q(rdata_c[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i6.GSR = "ENABLED";
    FD1P3AX rdata_i0_i5 (.D(n7958), .SP(n32444), .CK(debug_c_c), .Q(rdata_c[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i5.GSR = "ENABLED";
    FD1P3AX rdata_i0_i4 (.D(n7956), .SP(n32444), .CK(debug_c_c), .Q(rdata_c[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i4.GSR = "ENABLED";
    FD1P3AX rdata_i0_i3 (.D(n7954), .SP(n32444), .CK(debug_c_c), .Q(rdata_c[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i3.GSR = "ENABLED";
    FD1P3AX rdata_i0_i2 (.D(n7952), .SP(n32444), .CK(debug_c_c), .Q(rdata_c[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i2.GSR = "ENABLED";
    FD1P3AX rdata_i0_i1 (.D(n7950), .SP(n32444), .CK(debug_c_c), .Q(\rdata[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=27, LSE_RCOL=39, LSE_LLINE=60, LSE_RLINE=64 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam rdata_i0_i1.GSR = "ENABLED";
    LUT4 n30396_bdd_4_lut (.A(n32449), .B(state[4]), .C(bclk), .D(n32450), 
         .Z(n31419)) /* synthesis lut_function=(!((B (C (D))+!B !(C (D)))+!A)) */ ;
    defparam n30396_bdd_4_lut.init = 16'h2888;
    LUT4 i1_4_lut (.A(n11696), .B(rdata_c[2]), .C(n78[2]), .D(n13), 
         .Z(n7952)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i3699_4_lut (.A(n9396_c), .B(rdata_c[2]), .C(n11875), .D(n30516), 
         .Z(n78[2])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3699_4_lut.init = 16'hccca;
    LUT4 i1_4_lut_adj_26 (.A(n11696), .B(\rdata[1] ), .C(n31442), .D(n13), 
         .Z(n7950)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_26.init = 16'heca0;
    FD1S3IX drdy_51 (.D(n29148), .CK(debug_c_c), .CD(n34319), .Q(debug_c_7));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam drdy_51.GSR = "ENABLED";
    LUT4 i2927_3_lut_rep_399 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n32493)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2927_3_lut_rep_399.init = 16'h8080;
    LUT4 i2934_2_lut_rep_356_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(state[3]), .Z(n32450)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2934_2_lut_rep_356_4_lut.init = 16'h8000;
    LUT4 i21590_4_lut (.A(n183), .B(state[5]), .C(n1[3]), .D(n32), .Z(n29)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i21590_4_lut.init = 16'h3111;
    LUT4 i1_4_lut_adj_27 (.A(n11696), .B(rdata[0]), .C(n31427), .D(n13), 
         .Z(n7934)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_27.init = 16'heca0;
    LUT4 i2_3_lut (.A(state[0]), .B(state[4]), .C(state[5]), .Z(n11696)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i2_3_lut.init = 16'h0404;
    LUT4 i1_4_lut_adj_28 (.A(state[4]), .B(state[3]), .C(state[2]), .D(state[1]), 
         .Z(n32)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_28.init = 16'heaaa;
    LUT4 i2_3_lut_adj_29 (.A(state[0]), .B(state[5]), .C(state[4]), .Z(n13)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i2_3_lut_adj_29.init = 16'hefef;
    LUT4 i1_4_lut_4_lut (.A(state[5]), .B(n32432), .C(n9396_c), .D(debug_c_7), 
         .Z(n29148)) /* synthesis lut_function=(A ((D)+!B)+!A (B (D)+!B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_4_lut.init = 16'hfe22;
    LUT4 i1_4_lut_adj_30 (.A(state[5]), .B(state[2]), .C(n183), .D(n32), 
         .Z(n21)) /* synthesis lut_function=(!(A+!(B ((D)+!C)+!B !(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_30.init = 16'h4505;
    LUT4 i33_3_lut (.A(state[1]), .B(state[2]), .C(bclk), .Z(n17)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i33_3_lut.init = 16'hc6c6;
    LUT4 i2_4_lut (.A(bclk), .B(n4), .C(state[0]), .D(n32), .Z(n21_adj_7)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i2_4_lut.init = 16'h4840;
    LUT4 i38_4_lut (.A(n183), .B(n32450), .C(state[0]), .D(n4_adj_8), 
         .Z(n23)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (((D)+!C)+!B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i38_4_lut.init = 16'hf535;
    LUT4 i1_2_lut (.A(state[4]), .B(bclk), .Z(n4_adj_8)) /* synthesis lut_function=((B)+!A) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut.init = 16'hdddd;
    LUT4 i1_4_lut_adj_31 (.A(rdata[0]), .B(rx_data[0]), .C(n32409), .D(n19), 
         .Z(n7936)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_31.init = 16'heca0;
    LUT4 i4_4_lut (.A(n32495), .B(n32494), .C(state[5]), .D(state[0]), 
         .Z(n19)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i4_4_lut.init = 16'hffef;
    LUT4 i1_4_lut_adj_32 (.A(baud_reset), .B(n55), .C(n27961), .D(n56), 
         .Z(n2687)) /* synthesis lut_function=(A+!(B+((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_4_lut_adj_32.init = 16'haaba;
    LUT4 i1_2_lut_adj_33 (.A(state[1]), .B(bclk), .Z(n11875)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_33.init = 16'hbbbb;
    LUT4 i13_4_lut (.A(state[5]), .B(baud_reset), .C(n32432), .D(n9396_c), 
         .Z(n29398)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i13_4_lut.init = 16'hceca;
    LUT4 i1_2_lut_adj_34 (.A(state[1]), .B(bclk), .Z(n23288)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_34.init = 16'h8888;
    LUT4 i1_4_lut_adj_35 (.A(rdata_c[7]), .B(rx_data[7]), .C(n32409), 
         .D(n19), .Z(n7976)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_35.init = 16'heca0;
    LUT4 i1_4_lut_adj_36 (.A(rdata_c[6]), .B(rx_data[6]), .C(n32409), 
         .D(n19), .Z(n7974)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_36.init = 16'heca0;
    LUT4 i1_4_lut_adj_37 (.A(rdata_c[5]), .B(rx_data[5]), .C(n32409), 
         .D(n19), .Z(n7972)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_37.init = 16'heca0;
    LUT4 i1_4_lut_adj_38 (.A(rdata_c[4]), .B(rx_data[4]), .C(n32409), 
         .D(n19), .Z(n7970)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_38.init = 16'heca0;
    LUT4 i1_4_lut_adj_39 (.A(rdata_c[3]), .B(rx_data[3]), .C(n32409), 
         .D(n19), .Z(n7968)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_39.init = 16'heca0;
    LUT4 i1_4_lut_adj_40 (.A(rdata_c[2]), .B(rx_data[2]), .C(n32409), 
         .D(n19), .Z(n7966)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_40.init = 16'heca0;
    LUT4 i1_4_lut_adj_41 (.A(\rdata[1] ), .B(rx_data[1]), .C(n32409), 
         .D(n19), .Z(n7964)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_41.init = 16'heca0;
    LUT4 i1_4_lut_adj_42 (.A(n78[7]), .B(rdata_c[7]), .C(n11696), .D(n13), 
         .Z(n7962)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_42.init = 16'heca0;
    LUT4 i3689_4_lut (.A(rdata_c[7]), .B(n9396_c), .C(n23288), .D(n219), 
         .Z(n78[7])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3689_4_lut.init = 16'hcaaa;
    LUT4 i1_2_lut_adj_43 (.A(state[2]), .B(state[3]), .Z(n219)) /* synthesis lut_function=(A (B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_2_lut_adj_43.init = 16'h8888;
    LUT4 i1_4_lut_adj_44 (.A(n78[6]), .B(rdata_c[6]), .C(n11696), .D(n13), 
         .Z(n7960)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_44.init = 16'heca0;
    PFUMX i24897 (.BLUT(n31419), .ALUT(n31418), .C0(state[0]), .Z(n31420));
    LUT4 i3691_4_lut (.A(n9396_c), .B(rdata_c[6]), .C(n11875), .D(n219), 
         .Z(n78[6])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3691_4_lut.init = 16'hcacc;
    LUT4 i1_4_lut_adj_45 (.A(n78[5]), .B(rdata_c[5]), .C(n11696), .D(n13), 
         .Z(n7958)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_45.init = 16'heca0;
    LUT4 i3693_4_lut (.A(n9396_c), .B(rdata_c[5]), .C(state[1]), .D(n30483), 
         .Z(n78[5])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3693_4_lut.init = 16'hccac;
    LUT4 i1_3_lut (.A(state[2]), .B(state[3]), .C(bclk), .Z(n30483)) /* synthesis lut_function=(A+!(B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(29[9] 84[6])
    defparam i1_3_lut.init = 16'hbfbf;
    LUT4 i1_4_lut_adj_46 (.A(n78[4]), .B(rdata_c[4]), .C(n11696), .D(n13), 
         .Z(n7956)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_46.init = 16'heca0;
    LUT4 i3695_4_lut (.A(n9396_c), .B(rdata_c[4]), .C(state[1]), .D(n30483), 
         .Z(n78[4])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3695_4_lut.init = 16'hccca;
    LUT4 i1_4_lut_adj_47 (.A(n11696), .B(rdata_c[3]), .C(n78[3]), .D(n13), 
         .Z(n7954)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(39[6] 82[13])
    defparam i1_4_lut_adj_47.init = 16'heca0;
    LUT4 i3697_4_lut (.A(n9396_c), .B(rdata_c[3]), .C(n23288), .D(n30516), 
         .Z(n78[3])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(64[8] 68[12])
    defparam i3697_4_lut.init = 16'hccac;
    LUT4 i1_2_lut_adj_48 (.A(state[3]), .B(state[2]), .Z(n30516)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(67[10:27])
    defparam i1_2_lut_adj_48.init = 16'hbbbb;
    \ClockDividerP(factor=12)_U0  baud_gen (.bclk(bclk), .debug_c_c(debug_c_c), 
            .baud_reset(baud_reset), .n2687(n2687), .n55(n55), .n27961(n27961), 
            .n56(n56), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uart.v(25[28] 27[56])
    
endmodule
//
// Verilog Description of module \ClockDividerP(factor=12)_U0 
//

module \ClockDividerP(factor=12)_U0  (bclk, debug_c_c, baud_reset, n2687, 
            n55, n27961, n56, GND_net) /* synthesis syn_module_defined=1 */ ;
    output bclk;
    input debug_c_c;
    input baud_reset;
    input n2687;
    output n55;
    output n27961;
    output n56;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n7229;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(13[13:18])
    wire [31:0]n134;
    
    wire n52, n44, n35, n54, n48, n36, n46, n32, n50, n40, 
        n27537, n27536, n27535, n27534, n27533, n27532, n27531, 
        n27530, n27529, n27528, n27527, n27845, n27526, n27844, 
        n27843, n27525, n27842, n27841, n27524, n27840, n27839, 
        n27523, n27838, n27837, n27522, n27836, n27835, n27834, 
        n27833, n27832, n27831, n27830;
    
    FD1S3IX clk_o_14 (.D(n7229), .CK(debug_c_c), .CD(baud_reset), .Q(bclk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(15[9] 34[6])
    defparam clk_o_14.GSR = "ENABLED";
    FD1S3IX count_2180__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2687), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i0.GSR = "ENABLED";
    FD1S3IX count_2180__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2687), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i1.GSR = "ENABLED";
    FD1S3IX count_2180__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2687), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i2.GSR = "ENABLED";
    FD1S3IX count_2180__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2687), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i3.GSR = "ENABLED";
    FD1S3IX count_2180__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2687), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i4.GSR = "ENABLED";
    FD1S3IX count_2180__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2687), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i5.GSR = "ENABLED";
    FD1S3IX count_2180__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2687), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i6.GSR = "ENABLED";
    FD1S3IX count_2180__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2687), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i7.GSR = "ENABLED";
    FD1S3IX count_2180__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2687), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i8.GSR = "ENABLED";
    FD1S3IX count_2180__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2687), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i9.GSR = "ENABLED";
    FD1S3IX count_2180__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i10.GSR = "ENABLED";
    FD1S3IX count_2180__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i11.GSR = "ENABLED";
    FD1S3IX count_2180__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i12.GSR = "ENABLED";
    FD1S3IX count_2180__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i13.GSR = "ENABLED";
    FD1S3IX count_2180__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i14.GSR = "ENABLED";
    FD1S3IX count_2180__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i15.GSR = "ENABLED";
    FD1S3IX count_2180__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i16.GSR = "ENABLED";
    FD1S3IX count_2180__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i17.GSR = "ENABLED";
    FD1S3IX count_2180__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i18.GSR = "ENABLED";
    FD1S3IX count_2180__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i19.GSR = "ENABLED";
    FD1S3IX count_2180__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i20.GSR = "ENABLED";
    FD1S3IX count_2180__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i21.GSR = "ENABLED";
    FD1S3IX count_2180__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i22.GSR = "ENABLED";
    FD1S3IX count_2180__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i23.GSR = "ENABLED";
    FD1S3IX count_2180__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i24.GSR = "ENABLED";
    FD1S3IX count_2180__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i25.GSR = "ENABLED";
    FD1S3IX count_2180__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i26.GSR = "ENABLED";
    FD1S3IX count_2180__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i27.GSR = "ENABLED";
    FD1S3IX count_2180__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i28.GSR = "ENABLED";
    FD1S3IX count_2180__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i29.GSR = "ENABLED";
    FD1S3IX count_2180__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i30.GSR = "ENABLED";
    FD1S3IX count_2180__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2687), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180__i31.GSR = "ENABLED";
    LUT4 i26_4_lut (.A(count[30]), .B(n52), .C(n44), .D(count[14]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut (.A(count[1]), .B(count[3]), .C(count[0]), .Z(n27961)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i27_4_lut (.A(n35), .B(n54), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i23_4_lut (.A(count[12]), .B(n46), .C(n32), .D(count[18]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i15_3_lut (.A(count[15]), .B(count[24]), .C(count[31]), .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i17_4_lut (.A(count[16]), .B(count[10]), .C(count[9]), .D(count[17]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[20]), .B(count[5]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(count[13]), .B(count[22]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i25_4_lut (.A(count[7]), .B(n50), .C(n40), .D(count[11]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(count[4]), .B(count[6]), .C(count[8]), .D(count[29]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count[26]), .B(count[28]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i21_4_lut (.A(count[25]), .B(count[23]), .C(count[2]), .D(count[27]), 
         .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i11_2_lut (.A(count[19]), .B(count[21]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i11_2_lut.init = 16'heeee;
    CCU2D sub_1734_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27537), .S0(n7229));
    defparam sub_1734_add_2_cout.INIT0 = 16'h0000;
    defparam sub_1734_add_2_cout.INIT1 = 16'h0000;
    defparam sub_1734_add_2_cout.INJECT1_0 = "NO";
    defparam sub_1734_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27536), .COUT(n27537));
    defparam sub_1734_add_2_32.INIT0 = 16'h5555;
    defparam sub_1734_add_2_32.INIT1 = 16'h5555;
    defparam sub_1734_add_2_32.INJECT1_0 = "NO";
    defparam sub_1734_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27535), .COUT(n27536));
    defparam sub_1734_add_2_30.INIT0 = 16'h5555;
    defparam sub_1734_add_2_30.INIT1 = 16'h5555;
    defparam sub_1734_add_2_30.INJECT1_0 = "NO";
    defparam sub_1734_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27534), .COUT(n27535));
    defparam sub_1734_add_2_28.INIT0 = 16'h5555;
    defparam sub_1734_add_2_28.INIT1 = 16'h5555;
    defparam sub_1734_add_2_28.INJECT1_0 = "NO";
    defparam sub_1734_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27533), .COUT(n27534));
    defparam sub_1734_add_2_26.INIT0 = 16'h5555;
    defparam sub_1734_add_2_26.INIT1 = 16'h5555;
    defparam sub_1734_add_2_26.INJECT1_0 = "NO";
    defparam sub_1734_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27532), .COUT(n27533));
    defparam sub_1734_add_2_24.INIT0 = 16'h5555;
    defparam sub_1734_add_2_24.INIT1 = 16'h5555;
    defparam sub_1734_add_2_24.INJECT1_0 = "NO";
    defparam sub_1734_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27531), .COUT(n27532));
    defparam sub_1734_add_2_22.INIT0 = 16'h5555;
    defparam sub_1734_add_2_22.INIT1 = 16'h5555;
    defparam sub_1734_add_2_22.INJECT1_0 = "NO";
    defparam sub_1734_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27530), .COUT(n27531));
    defparam sub_1734_add_2_20.INIT0 = 16'h5555;
    defparam sub_1734_add_2_20.INIT1 = 16'h5555;
    defparam sub_1734_add_2_20.INJECT1_0 = "NO";
    defparam sub_1734_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27529), .COUT(n27530));
    defparam sub_1734_add_2_18.INIT0 = 16'h5555;
    defparam sub_1734_add_2_18.INIT1 = 16'h5555;
    defparam sub_1734_add_2_18.INJECT1_0 = "NO";
    defparam sub_1734_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27528), .COUT(n27529));
    defparam sub_1734_add_2_16.INIT0 = 16'h5555;
    defparam sub_1734_add_2_16.INIT1 = 16'h5555;
    defparam sub_1734_add_2_16.INJECT1_0 = "NO";
    defparam sub_1734_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27527), .COUT(n27528));
    defparam sub_1734_add_2_14.INIT0 = 16'h5555;
    defparam sub_1734_add_2_14.INIT1 = 16'h5555;
    defparam sub_1734_add_2_14.INJECT1_0 = "NO";
    defparam sub_1734_add_2_14.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27845), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_33.INIT1 = 16'h0000;
    defparam count_2180_add_4_33.INJECT1_0 = "NO";
    defparam count_2180_add_4_33.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27526), .COUT(n27527));
    defparam sub_1734_add_2_12.INIT0 = 16'h5555;
    defparam sub_1734_add_2_12.INIT1 = 16'h5555;
    defparam sub_1734_add_2_12.INJECT1_0 = "NO";
    defparam sub_1734_add_2_12.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27844), .COUT(n27845), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_31.INJECT1_0 = "NO";
    defparam count_2180_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27843), .COUT(n27844), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_29.INJECT1_0 = "NO";
    defparam count_2180_add_4_29.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27525), .COUT(n27526));
    defparam sub_1734_add_2_10.INIT0 = 16'h5555;
    defparam sub_1734_add_2_10.INIT1 = 16'h5555;
    defparam sub_1734_add_2_10.INJECT1_0 = "NO";
    defparam sub_1734_add_2_10.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27842), .COUT(n27843), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_27.INJECT1_0 = "NO";
    defparam count_2180_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27841), .COUT(n27842), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_25.INJECT1_0 = "NO";
    defparam count_2180_add_4_25.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27524), .COUT(n27525));
    defparam sub_1734_add_2_8.INIT0 = 16'h5555;
    defparam sub_1734_add_2_8.INIT1 = 16'h5555;
    defparam sub_1734_add_2_8.INJECT1_0 = "NO";
    defparam sub_1734_add_2_8.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27840), .COUT(n27841), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_23.INJECT1_0 = "NO";
    defparam count_2180_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27839), .COUT(n27840), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_21.INJECT1_0 = "NO";
    defparam count_2180_add_4_21.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27523), .COUT(n27524));
    defparam sub_1734_add_2_6.INIT0 = 16'h5555;
    defparam sub_1734_add_2_6.INIT1 = 16'h5555;
    defparam sub_1734_add_2_6.INJECT1_0 = "NO";
    defparam sub_1734_add_2_6.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27838), .COUT(n27839), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_19.INJECT1_0 = "NO";
    defparam count_2180_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27837), .COUT(n27838), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_17.INJECT1_0 = "NO";
    defparam count_2180_add_4_17.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27522), .COUT(n27523));
    defparam sub_1734_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_1734_add_2_4.INIT1 = 16'h5555;
    defparam sub_1734_add_2_4.INJECT1_0 = "NO";
    defparam sub_1734_add_2_4.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27836), .COUT(n27837), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_15.INJECT1_0 = "NO";
    defparam count_2180_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27835), .COUT(n27836), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_13.INJECT1_0 = "NO";
    defparam count_2180_add_4_13.INJECT1_1 = "NO";
    CCU2D sub_1734_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27522));
    defparam sub_1734_add_2_2.INIT0 = 16'h0000;
    defparam sub_1734_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_1734_add_2_2.INJECT1_0 = "NO";
    defparam sub_1734_add_2_2.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27834), .COUT(n27835), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_11.INJECT1_0 = "NO";
    defparam count_2180_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27833), .COUT(n27834), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_9.INJECT1_0 = "NO";
    defparam count_2180_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27832), .COUT(n27833), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_7.INJECT1_0 = "NO";
    defparam count_2180_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27831), .COUT(n27832), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_5.INJECT1_0 = "NO";
    defparam count_2180_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27830), .COUT(n27831), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2180_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2180_add_4_3.INJECT1_0 = "NO";
    defparam count_2180_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2180_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27830), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(32[16:25])
    defparam count_2180_add_4_1.INIT0 = 16'hF000;
    defparam count_2180_add_4_1.INIT1 = 16'h0555;
    defparam count_2180_add_4_1.INJECT1_0 = "NO";
    defparam count_2180_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \ArmPeripheral(axis_haddr=8'b0) 
//

module \ArmPeripheral(axis_haddr=8'b0)  (\register_addr[0] , debug_c_c, 
            n34324, n3451, n32401, prev_select, \register_addr[5] , 
            n34317, n32343, n34321, limit_c_0, n32481, n32480, n32460, 
            n302, \register_addr[1] , n32504, n30726, n32422, \read_size[0] , 
            n11966, n34322, Stepper_X_M0_c_0, n579, n34323, \steps_reg[7] , 
            read_value, \databus[31] , n34325, \databus[30] , \databus[29] , 
            \databus[26] , \databus[13] , \databus[11] , \databus[10] , 
            \databus[9] , \databus[7] , \databus[6] , \databus[5] , 
            n608, n610, \control_reg[7] , Stepper_X_En_c, n34326, 
            Stepper_X_Dir_c, \databus[3] , Stepper_X_M2_c_2, Stepper_X_M1_c_1, 
            \databus[1] , \read_size[2] , n32433, \register_addr[4] , 
            \register_addr[3] , n11753, n30310, n30313, n11645, n34320, 
            GND_net, n224, n21, n30423, n32365, n12434, \register_addr[6] , 
            \register_addr[7] , n32448, n32503, n20268, n28356, \databus[8] , 
            \databus[12] , \databus[14] , \databus[15] , n32455, n32442, 
            n32369, rw, n32350, \databus[16] , \databus[17] , \databus[18] , 
            \databus[19] , \databus[20] , \databus[21] , \databus[22] , 
            \databus[23] , n32354, \databus[24] , \databus[25] , \databus[27] , 
            \databus[28] , VCC_net, Stepper_X_nFault_c, n28332, n32379, 
            n30401, n8048, n13, Stepper_X_Step_c) /* synthesis syn_module_defined=1 */ ;
    input \register_addr[0] ;
    input debug_c_c;
    input n34324;
    input [31:0]n3451;
    input n32401;
    output prev_select;
    input \register_addr[5] ;
    input n34317;
    output n32343;
    input n34321;
    input limit_c_0;
    output n32481;
    input n32480;
    input n32460;
    output n302;
    input \register_addr[1] ;
    input n32504;
    output n30726;
    output n32422;
    output \read_size[0] ;
    input n11966;
    input n34322;
    output Stepper_X_M0_c_0;
    input n579;
    input n34323;
    output \steps_reg[7] ;
    output [31:0]read_value;
    input \databus[31] ;
    input n34325;
    input \databus[30] ;
    input \databus[29] ;
    input \databus[26] ;
    input \databus[13] ;
    input \databus[11] ;
    input \databus[10] ;
    input \databus[9] ;
    input \databus[7] ;
    input \databus[6] ;
    input \databus[5] ;
    input n608;
    input n610;
    output \control_reg[7] ;
    output Stepper_X_En_c;
    input n34326;
    output Stepper_X_Dir_c;
    input \databus[3] ;
    output Stepper_X_M2_c_2;
    output Stepper_X_M1_c_1;
    input \databus[1] ;
    output \read_size[2] ;
    input n32433;
    input \register_addr[4] ;
    input \register_addr[3] ;
    input n11753;
    output n30310;
    input n30313;
    output n11645;
    input n34320;
    input GND_net;
    output [31:0]n224;
    input n21;
    input n30423;
    input n32365;
    output n12434;
    input \register_addr[6] ;
    input \register_addr[7] ;
    output n32448;
    input n32503;
    input n20268;
    output n28356;
    input \databus[8] ;
    input \databus[12] ;
    input \databus[14] ;
    input \databus[15] ;
    input n32455;
    input n32442;
    input n32369;
    input rw;
    input n32350;
    input \databus[16] ;
    input \databus[17] ;
    input \databus[18] ;
    input \databus[19] ;
    input \databus[20] ;
    input \databus[21] ;
    input \databus[22] ;
    input \databus[23] ;
    input n32354;
    input \databus[24] ;
    input \databus[25] ;
    input \databus[27] ;
    input \databus[28] ;
    input VCC_net;
    input Stepper_X_nFault_c;
    output n28332;
    input n32379;
    input n30401;
    output n8048;
    input n13;
    output Stepper_X_Step_c;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n30863, n30864, n30865;
    wire [31:0]steps_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(28[13:22])
    
    wire n182, n30169, n12540, prev_step_clk, step_clk, limit_latched, 
        prev_limit_latched;
    wire [31:0]div_factor_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(27[13:27])
    
    wire n12480, n30314, n30318, n30316, n30317, n30315, n30319, 
        n30329, n30328, n30330, n30331, n30332, n30333, n30334, 
        n30335, n30336, n30337, n32342, n32349, n9614;
    wire [7:0]control_reg;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(26[12:23])
    
    wire n1, n2, n32465, n17324, int_step, n12, n32362, n27746, 
        n27747, n27745, n27744, n27743, n27742, n1_adj_1, n2_adj_2;
    wire [31:0]n5188;
    
    wire n1_adj_3, n2_adj_4, n1_adj_5, n2_adj_6, n30856, n30853, 
        n30327, n30326, n30325, n30324, n30323, n30322, n30321, 
        fault_latched, n30854, n30855, n30851, n30852, n30320, n49, 
        n62, n58, n50, n41, n60, n54, n42, n52, n38, n56, 
        n46, n27757, n27756, n27755, n27754, n27753, n27752, n27751, 
        n27750, n27749, n27748;
    
    PFUMX i24506 (.BLUT(n30863), .ALUT(n30864), .C0(\register_addr[0] ), 
          .Z(n30865));
    FD1S3IX steps_reg__i19 (.D(n3451[19]), .CK(debug_c_c), .CD(n34324), 
            .Q(steps_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i19.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_249_3_lut_4_lut (.A(n32401), .B(prev_select), .C(\register_addr[5] ), 
         .D(n34317), .Z(n32343)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(82[9:30])
    defparam i1_2_lut_rep_249_3_lut_4_lut.init = 16'h0002;
    FD1S3IX steps_reg__i18 (.D(n3451[18]), .CK(debug_c_c), .CD(n34321), 
            .Q(steps_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i18.GSR = "ENABLED";
    LUT4 i118_1_lut (.A(limit_c_0), .Z(n182)) /* synthesis lut_function=(!(A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(62[21:28])
    defparam i118_1_lut.init = 16'h5555;
    FD1S3IX steps_reg__i17 (.D(n3451[17]), .CK(debug_c_c), .CD(n34321), 
            .Q(steps_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i17.GSR = "ENABLED";
    FD1S3IX steps_reg__i16 (.D(n3451[16]), .CK(debug_c_c), .CD(n34321), 
            .Q(steps_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i16.GSR = "ENABLED";
    FD1S3IX steps_reg__i0 (.D(n3451[0]), .CK(debug_c_c), .CD(n34321), 
            .Q(steps_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i0.GSR = "ENABLED";
    FD1S3IX steps_reg__i15 (.D(n3451[15]), .CK(debug_c_c), .CD(n34321), 
            .Q(steps_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i15.GSR = "ENABLED";
    FD1S3IX steps_reg__i14 (.D(n3451[14]), .CK(debug_c_c), .CD(n34321), 
            .Q(steps_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i14.GSR = "ENABLED";
    LUT4 equal_138_i16_1_lut_2_lut_3_lut_4_lut (.A(n32481), .B(n32480), 
         .C(n32460), .D(\register_addr[0] ), .Z(n302)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam equal_138_i16_1_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32481), .B(n32480), .C(\register_addr[1] ), 
         .D(n32504), .Z(n30169)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i24805_2_lut_3_lut_4_lut (.A(n32481), .B(n32480), .C(\register_addr[1] ), 
         .D(n32504), .Z(n30726)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i24805_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 equal_138_i15_2_lut_rep_328_3_lut_4_lut (.A(n32481), .B(n32480), 
         .C(n32460), .D(\register_addr[0] ), .Z(n32422)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam equal_138_i15_2_lut_rep_328_3_lut_4_lut.init = 16'hfffe;
    FD1P3AX read_size__i1 (.D(n30726), .SP(n11966), .CK(debug_c_c), .Q(\read_size[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i1.GSR = "ENABLED";
    FD1S3IX steps_reg__i13 (.D(n3451[13]), .CK(debug_c_c), .CD(n34322), 
            .Q(steps_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i13.GSR = "ENABLED";
    FD1S3IX steps_reg__i12 (.D(n3451[12]), .CK(debug_c_c), .CD(n34322), 
            .Q(steps_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i12.GSR = "ENABLED";
    FD1P3AX control_reg_i1 (.D(n579), .SP(n12540), .CK(debug_c_c), .Q(Stepper_X_M0_c_0)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i1.GSR = "ENABLED";
    FD1S3AX prev_step_clk_175 (.D(step_clk), .CK(debug_c_c), .Q(prev_step_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_step_clk_175.GSR = "ENABLED";
    FD1S3AX limit_latched_176 (.D(n182), .CK(debug_c_c), .Q(limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam limit_latched_176.GSR = "ENABLED";
    FD1S3AX prev_limit_latched_177 (.D(limit_latched), .CK(debug_c_c), .Q(prev_limit_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_limit_latched_177.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i0 (.D(n579), .SP(n12480), .CK(debug_c_c), 
            .Q(div_factor_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i0.GSR = "ENABLED";
    FD1S3IX steps_reg__i11 (.D(n3451[11]), .CK(debug_c_c), .CD(n34322), 
            .Q(steps_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i11.GSR = "ENABLED";
    FD1S3AX prev_select_174 (.D(n32401), .CK(debug_c_c), .Q(prev_select)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam prev_select_174.GSR = "ENABLED";
    FD1S3IX steps_reg__i10 (.D(n3451[10]), .CK(debug_c_c), .CD(n34322), 
            .Q(steps_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i10.GSR = "ENABLED";
    FD1S3IX steps_reg__i9 (.D(n3451[9]), .CK(debug_c_c), .CD(n34322), 
            .Q(steps_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i9.GSR = "ENABLED";
    FD1S3IX steps_reg__i8 (.D(n3451[8]), .CK(debug_c_c), .CD(n34323), 
            .Q(steps_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i8.GSR = "ENABLED";
    FD1S3IX steps_reg__i7 (.D(n3451[7]), .CK(debug_c_c), .CD(n34323), 
            .Q(\steps_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i7.GSR = "ENABLED";
    FD1S3IX steps_reg__i6 (.D(n3451[6]), .CK(debug_c_c), .CD(n34323), 
            .Q(steps_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i6.GSR = "ENABLED";
    FD1S3IX steps_reg__i5 (.D(n3451[5]), .CK(debug_c_c), .CD(n34323), 
            .Q(steps_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i5.GSR = "ENABLED";
    FD1S3IX steps_reg__i4 (.D(n3451[4]), .CK(debug_c_c), .CD(n34323), 
            .Q(steps_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i4.GSR = "ENABLED";
    FD1S3IX steps_reg__i3 (.D(n3451[3]), .CK(debug_c_c), .CD(n34323), 
            .Q(steps_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i3.GSR = "ENABLED";
    FD1S3IX steps_reg__i2 (.D(n3451[2]), .CK(debug_c_c), .CD(n34323), 
            .Q(steps_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i1 (.D(n3451[1]), .CK(debug_c_c), .CD(n34323), 
            .Q(steps_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i1.GSR = "ENABLED";
    FD1P3AX read_value__i16 (.D(n30314), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i16.GSR = "ENABLED";
    FD1P3AX read_value__i17 (.D(n30318), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i17.GSR = "ENABLED";
    FD1P3AX read_value__i18 (.D(n30316), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i18.GSR = "ENABLED";
    FD1P3AX read_value__i19 (.D(n30317), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i19.GSR = "ENABLED";
    FD1P3AX read_value__i20 (.D(n30315), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i20.GSR = "ENABLED";
    FD1P3AX read_value__i21 (.D(n30319), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i21.GSR = "ENABLED";
    FD1P3AX read_value__i22 (.D(n30329), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i22.GSR = "ENABLED";
    FD1P3AX read_value__i23 (.D(n30328), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i23.GSR = "ENABLED";
    FD1P3AX read_value__i24 (.D(n30330), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i24.GSR = "ENABLED";
    FD1P3AX read_value__i25 (.D(n30331), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i25.GSR = "ENABLED";
    FD1P3AX read_value__i26 (.D(n30332), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i26.GSR = "ENABLED";
    FD1P3AX read_value__i27 (.D(n30333), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i27.GSR = "ENABLED";
    FD1P3AX read_value__i28 (.D(n30334), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i28.GSR = "ENABLED";
    FD1P3AX read_value__i29 (.D(n30335), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i29.GSR = "ENABLED";
    FD1P3AX read_value__i30 (.D(n30336), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i30.GSR = "ENABLED";
    FD1P3AX read_value__i31 (.D(n30337), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i31 (.D(\databus[31] ), .SP(n32342), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i31.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i30 (.D(\databus[30] ), .SP(n32342), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i30.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i29 (.D(\databus[29] ), .SP(n32342), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i29.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i26 (.D(\databus[26] ), .SP(n32342), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i26.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i13 (.D(\databus[13] ), .SP(n32342), .PD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i13.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i11 (.D(\databus[11] ), .SP(n32342), .PD(n34324), 
            .CK(debug_c_c), .Q(div_factor_reg[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i11.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i10 (.D(\databus[10] ), .SP(n32342), .PD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i10.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i9 (.D(\databus[9] ), .SP(n32342), .PD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i9.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i7 (.D(\databus[7] ), .SP(n32342), .PD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i7.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i6 (.D(\databus[6] ), .SP(n32342), .PD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i6.GSR = "ENABLED";
    FD1P3JX div_factor_reg_i5 (.D(\databus[5] ), .SP(n32342), .PD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i5.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i4 (.D(n608), .SP(n12480), .CK(debug_c_c), 
            .Q(div_factor_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i4.GSR = "ENABLED";
    FD1P3AX div_factor_reg_i2 (.D(n610), .SP(n12480), .CK(debug_c_c), 
            .Q(div_factor_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i2.GSR = "ENABLED";
    FD1P3IX control_reg_i8 (.D(\databus[7] ), .SP(n32349), .CD(n9614), 
            .CK(debug_c_c), .Q(\control_reg[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i8.GSR = "ENABLED";
    FD1P3JX control_reg_i7 (.D(\databus[6] ), .SP(n32349), .PD(n34326), 
            .CK(debug_c_c), .Q(Stepper_X_En_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i7.GSR = "ENABLED";
    FD1P3JX control_reg_i6 (.D(\databus[5] ), .SP(n32349), .PD(n34326), 
            .CK(debug_c_c), .Q(Stepper_X_Dir_c)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i6.GSR = "ENABLED";
    FD1P3AX control_reg_i5 (.D(n608), .SP(n12540), .CK(debug_c_c), .Q(control_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i5.GSR = "ENABLED";
    FD1P3JX control_reg_i4 (.D(\databus[3] ), .SP(n32349), .PD(n34326), 
            .CK(debug_c_c), .Q(control_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i4.GSR = "ENABLED";
    FD1P3AX control_reg_i3 (.D(n610), .SP(n12540), .CK(debug_c_c), .Q(Stepper_X_M2_c_2)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i3.GSR = "ENABLED";
    FD1P3JX control_reg_i2 (.D(\databus[1] ), .SP(n32349), .PD(n34326), 
            .CK(debug_c_c), .Q(Stepper_X_M1_c_1)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam control_reg_i2.GSR = "ENABLED";
    FD1P3AX read_size__i2 (.D(n30169), .SP(n11966), .CK(debug_c_c), .Q(\read_size[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_size__i2.GSR = "ENABLED";
    FD1S3IX steps_reg__i31 (.D(n3451[31]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[31])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i31.GSR = "ENABLED";
    LUT4 i14201_2_lut (.A(Stepper_X_En_c), .B(\register_addr[0] ), .Z(n1)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14201_2_lut.init = 16'h2222;
    LUT4 mux_1600_Mux_6_i2_3_lut (.A(div_factor_reg[6]), .B(steps_reg[6]), 
         .C(\register_addr[0] ), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1600_Mux_6_i2_3_lut.init = 16'hcaca;
    FD1S3IX steps_reg__i30 (.D(n3451[30]), .CK(debug_c_c), .CD(n34326), 
            .Q(steps_reg[30])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i30.GSR = "ENABLED";
    FD1S3IX steps_reg__i29 (.D(n3451[29]), .CK(debug_c_c), .CD(n32433), 
            .Q(steps_reg[29])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i29.GSR = "ENABLED";
    FD1S3IX steps_reg__i28 (.D(n3451[28]), .CK(debug_c_c), .CD(n32433), 
            .Q(steps_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i28.GSR = "ENABLED";
    FD1S3IX steps_reg__i27 (.D(n3451[27]), .CK(debug_c_c), .CD(n32433), 
            .Q(steps_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i27.GSR = "ENABLED";
    FD1S3IX steps_reg__i26 (.D(n3451[26]), .CK(debug_c_c), .CD(n32433), 
            .Q(steps_reg[26])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i26.GSR = "ENABLED";
    FD1S3IX steps_reg__i25 (.D(n3451[25]), .CK(debug_c_c), .CD(n32433), 
            .Q(steps_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i25.GSR = "ENABLED";
    FD1S3IX steps_reg__i24 (.D(n3451[24]), .CK(debug_c_c), .CD(n32433), 
            .Q(steps_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i24.GSR = "ENABLED";
    FD1S3IX steps_reg__i23 (.D(n3451[23]), .CK(debug_c_c), .CD(n32433), 
            .Q(steps_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i23.GSR = "ENABLED";
    FD1S3IX steps_reg__i22 (.D(n3451[22]), .CK(debug_c_c), .CD(n32433), 
            .Q(steps_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i22.GSR = "ENABLED";
    FD1S3IX steps_reg__i21 (.D(n3451[21]), .CK(debug_c_c), .CD(n32433), 
            .Q(steps_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i21.GSR = "ENABLED";
    FD1S3IX steps_reg__i20 (.D(n3451[20]), .CK(debug_c_c), .CD(n32433), 
            .Q(steps_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam steps_reg__i20.GSR = "ENABLED";
    LUT4 i14218_2_lut_rep_371 (.A(\register_addr[4] ), .B(\register_addr[3] ), 
         .Z(n32465)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14218_2_lut_rep_371.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(\register_addr[4] ), .B(\register_addr[3] ), 
         .C(n11753), .Z(n30310)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_4_lut (.A(div_factor_reg[24]), .B(n30313), .C(steps_reg[24]), 
         .D(\register_addr[0] ), .Z(n30330)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_1 (.A(div_factor_reg[25]), .B(n30313), .C(steps_reg[25]), 
         .D(\register_addr[0] ), .Z(n30331)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_1.init = 16'hc088;
    LUT4 i1_4_lut_adj_2 (.A(div_factor_reg[26]), .B(n30313), .C(steps_reg[26]), 
         .D(\register_addr[0] ), .Z(n30332)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_2.init = 16'hc088;
    LUT4 i1_2_lut (.A(\register_addr[1] ), .B(\register_addr[0] ), .Z(n11645)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_3 (.A(div_factor_reg[27]), .B(n30313), .C(steps_reg[27]), 
         .D(\register_addr[0] ), .Z(n30333)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_3.init = 16'hc088;
    LUT4 i1_4_lut_adj_4 (.A(div_factor_reg[28]), .B(n30313), .C(steps_reg[28]), 
         .D(\register_addr[0] ), .Z(n30334)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_4.init = 16'hc088;
    LUT4 i1_4_lut_adj_5 (.A(div_factor_reg[29]), .B(n30313), .C(steps_reg[29]), 
         .D(\register_addr[0] ), .Z(n30335)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_5.init = 16'hc088;
    LUT4 i1_4_lut_adj_6 (.A(div_factor_reg[30]), .B(n30313), .C(steps_reg[30]), 
         .D(\register_addr[0] ), .Z(n30336)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_6.init = 16'hc088;
    LUT4 i1_4_lut_adj_7 (.A(div_factor_reg[31]), .B(n30313), .C(steps_reg[31]), 
         .D(\register_addr[0] ), .Z(n30337)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_7.init = 16'hc088;
    LUT4 i11573_3_lut (.A(\control_reg[7] ), .B(div_factor_reg[7]), .C(\register_addr[1] ), 
         .Z(n17324)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i11573_3_lut.init = 16'hcaca;
    LUT4 i3853_3_lut (.A(prev_limit_latched), .B(n34320), .C(limit_latched), 
         .Z(n9614)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(73[5] 127[8])
    defparam i3853_3_lut.init = 16'hdcdc;
    FD1P3AX int_step_182 (.D(n32362), .SP(n12), .CK(debug_c_c), .Q(int_step));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam int_step_182.GSR = "ENABLED";
    CCU2D sub_125_add_2_11 (.A0(steps_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27746), .COUT(n27747), .S0(n224[9]), .S1(n224[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_11.INIT0 = 16'h5555;
    defparam sub_125_add_2_11.INIT1 = 16'h5555;
    defparam sub_125_add_2_11.INJECT1_0 = "NO";
    defparam sub_125_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_9 (.A0(\steps_reg[7] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27745), .COUT(n27746), .S0(n224[7]), .S1(n224[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_9.INIT0 = 16'h5555;
    defparam sub_125_add_2_9.INIT1 = 16'h5555;
    defparam sub_125_add_2_9.INJECT1_0 = "NO";
    defparam sub_125_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_7 (.A0(steps_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27744), .COUT(n27745), .S0(n224[5]), .S1(n224[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_7.INIT0 = 16'h5555;
    defparam sub_125_add_2_7.INIT1 = 16'h5555;
    defparam sub_125_add_2_7.INJECT1_0 = "NO";
    defparam sub_125_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_5 (.A0(steps_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27743), .COUT(n27744), .S0(n224[3]), .S1(n224[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_5.INIT0 = 16'h5555;
    defparam sub_125_add_2_5.INIT1 = 16'h5555;
    defparam sub_125_add_2_5.INJECT1_0 = "NO";
    defparam sub_125_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_3 (.A0(steps_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27742), .COUT(n27743), .S0(n224[1]), .S1(n224[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_3.INIT0 = 16'h5555;
    defparam sub_125_add_2_3.INIT1 = 16'h5555;
    defparam sub_125_add_2_3.INJECT1_0 = "NO";
    defparam sub_125_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(steps_reg[0]), .B1(step_clk), .C1(n21), .D1(prev_step_clk), 
          .COUT(n27742), .S1(n224[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_1.INIT0 = 16'h0000;
    defparam sub_125_add_2_1.INIT1 = 16'h5595;
    defparam sub_125_add_2_1.INJECT1_0 = "NO";
    defparam sub_125_add_2_1.INJECT1_1 = "NO";
    PFUMX mux_1600_Mux_3_i3 (.BLUT(n1_adj_1), .ALUT(n2_adj_2), .C0(\register_addr[1] ), 
          .Z(n5188[3]));
    PFUMX mux_1600_Mux_4_i3 (.BLUT(n1_adj_3), .ALUT(n2_adj_4), .C0(\register_addr[1] ), 
          .Z(n5188[4]));
    PFUMX mux_1600_Mux_5_i3 (.BLUT(n1_adj_5), .ALUT(n2_adj_6), .C0(\register_addr[1] ), 
          .Z(n5188[5]));
    LUT4 i1_2_lut_4_lut (.A(n30423), .B(\register_addr[4] ), .C(n32365), 
         .D(n34320), .Z(n12434)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_2_lut_4_lut.init = 16'hff80;
    LUT4 equal_138_i13_2_lut_rep_387 (.A(\register_addr[6] ), .B(\register_addr[7] ), 
         .Z(n32481)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam equal_138_i13_2_lut_rep_387.init = 16'heeee;
    LUT4 i1_2_lut_rep_354_3_lut_4_lut (.A(\register_addr[6] ), .B(\register_addr[7] ), 
         .C(\register_addr[5] ), .D(\register_addr[4] ), .Z(n32448)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i1_2_lut_rep_354_3_lut_4_lut.init = 16'hfffe;
    LUT4 i24748_4_lut (.A(n32503), .B(n20268), .C(\register_addr[5] ), 
         .D(n32465), .Z(n28356)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i24748_4_lut.init = 16'h0001;
    FD1P3IX div_factor_reg_i1 (.D(\databus[1] ), .SP(n12480), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i1.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i3 (.D(\databus[3] ), .SP(n12480), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i3.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_8 (.A(div_factor_reg[16]), .B(n30313), .C(steps_reg[16]), 
         .D(\register_addr[0] ), .Z(n30314)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i1_4_lut_adj_8.init = 16'hc088;
    FD1P3IX div_factor_reg_i8 (.D(\databus[8] ), .SP(n12480), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i8.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i12 (.D(\databus[12] ), .SP(n12480), .CD(n34324), 
            .CK(debug_c_c), .Q(div_factor_reg[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i12.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i14 (.D(\databus[14] ), .SP(n12480), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i14.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_9 (.A(div_factor_reg[17]), .B(n30313), .C(steps_reg[17]), 
         .D(\register_addr[0] ), .Z(n30318)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_9.init = 16'hc088;
    FD1P3IX div_factor_reg_i15 (.D(\databus[15] ), .SP(n12480), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i15.GSR = "ENABLED";
    LUT4 i24726_3_lut_rep_255_4_lut_4_lut (.A(n32455), .B(n32442), .C(n32369), 
         .D(rw), .Z(n32349)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i24726_3_lut_rep_255_4_lut_4_lut.init = 16'h0010;
    LUT4 i24716_2_lut_4_lut_4_lut (.A(n32455), .B(n34320), .C(n32350), 
         .D(n32442), .Z(n12540)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(114[11:28])
    defparam i24716_2_lut_4_lut_4_lut.init = 16'hccdc;
    FD1P3IX div_factor_reg_i16 (.D(\databus[16] ), .SP(n12480), .CD(n34324), 
            .CK(debug_c_c), .Q(div_factor_reg[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i16.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i17 (.D(\databus[17] ), .SP(n12480), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i17.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i18 (.D(\databus[18] ), .SP(n12480), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i18.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i19 (.D(\databus[19] ), .SP(n12480), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i19.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i20 (.D(\databus[20] ), .SP(n12480), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i20.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i21 (.D(\databus[21] ), .SP(n12480), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[21])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i21.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i22 (.D(\databus[22] ), .SP(n12480), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[22])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i22.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i23 (.D(\databus[23] ), .SP(n12480), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[23])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i23.GSR = "ENABLED";
    FD1P3IX read_value__i1 (.D(n30856), .SP(n11966), .CD(n32354), .CK(debug_c_c), 
            .Q(read_value[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i1.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_10 (.A(div_factor_reg[18]), .B(n30313), .C(steps_reg[18]), 
         .D(\register_addr[0] ), .Z(n30316)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_10.init = 16'hc088;
    LUT4 i1_4_lut_adj_11 (.A(div_factor_reg[19]), .B(n30313), .C(steps_reg[19]), 
         .D(\register_addr[0] ), .Z(n30317)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_11.init = 16'hc088;
    FD1P3IX read_value__i2 (.D(n30853), .SP(n11966), .CD(n32354), .CK(debug_c_c), 
            .Q(read_value[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i2.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut_adj_12 (.A(n30423), .B(\register_addr[4] ), .C(n32343), 
         .D(n34320), .Z(n12480)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;
    defparam i1_2_lut_4_lut_adj_12.init = 16'hff20;
    FD1P3IX read_value__i3 (.D(n5188[3]), .SP(n11966), .CD(n32354), .CK(debug_c_c), 
            .Q(read_value[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i3.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i24 (.D(\databus[24] ), .SP(n12480), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[24])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i24.GSR = "ENABLED";
    FD1P3IX read_value__i4 (.D(n5188[4]), .SP(n11966), .CD(n32354), .CK(debug_c_c), 
            .Q(read_value[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i4.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i25 (.D(\databus[25] ), .SP(n12480), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[25])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i25.GSR = "ENABLED";
    FD1P3IX read_value__i5 (.D(n5188[5]), .SP(n11966), .CD(n32354), .CK(debug_c_c), 
            .Q(read_value[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i5.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i27 (.D(\databus[27] ), .SP(n12480), .CD(n34321), 
            .CK(debug_c_c), .Q(div_factor_reg[27])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i27.GSR = "ENABLED";
    FD1P3IX read_value__i6 (.D(n5188[6]), .SP(n11966), .CD(n32354), .CK(debug_c_c), 
            .Q(read_value[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i6.GSR = "ENABLED";
    FD1P3IX div_factor_reg_i28 (.D(\databus[28] ), .SP(n12480), .CD(n34325), 
            .CK(debug_c_c), .Q(div_factor_reg[28])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam div_factor_reg_i28.GSR = "ENABLED";
    FD1P3IX read_value__i7 (.D(n5188[7]), .SP(n11966), .CD(n32354), .CK(debug_c_c), 
            .Q(read_value[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i7.GSR = "ENABLED";
    FD1P3AX read_value__i8 (.D(n30327), .SP(n11966), .CK(debug_c_c), .Q(read_value[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i8.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_13 (.A(div_factor_reg[20]), .B(n30313), .C(steps_reg[20]), 
         .D(\register_addr[0] ), .Z(n30315)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_13.init = 16'hc088;
    LUT4 i1_4_lut_adj_14 (.A(div_factor_reg[21]), .B(n30313), .C(steps_reg[21]), 
         .D(\register_addr[0] ), .Z(n30319)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_14.init = 16'hc088;
    FD1P3AX read_value__i9 (.D(n30326), .SP(n11966), .CK(debug_c_c), .Q(read_value[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i9.GSR = "ENABLED";
    FD1P3AX read_value__i10 (.D(n30325), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i10.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_15 (.A(div_factor_reg[22]), .B(n30313), .C(steps_reg[22]), 
         .D(\register_addr[0] ), .Z(n30329)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_15.init = 16'hc088;
    LUT4 i1_4_lut_adj_16 (.A(div_factor_reg[23]), .B(n30313), .C(steps_reg[23]), 
         .D(\register_addr[0] ), .Z(n30328)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_16.init = 16'hc088;
    LUT4 i2_3_lut_rep_248_4_lut (.A(\register_addr[5] ), .B(n32350), .C(\register_addr[4] ), 
         .D(n30423), .Z(n32342)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_rep_248_4_lut.init = 16'h0400;
    LUT4 i14204_2_lut (.A(control_reg[3]), .B(\register_addr[0] ), .Z(n1_adj_1)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14204_2_lut.init = 16'h2222;
    LUT4 mux_1600_Mux_3_i2_3_lut (.A(div_factor_reg[3]), .B(steps_reg[3]), 
         .C(\register_addr[0] ), .Z(n2_adj_2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1600_Mux_3_i2_3_lut.init = 16'hcaca;
    LUT4 i14203_2_lut (.A(control_reg[4]), .B(\register_addr[0] ), .Z(n1_adj_3)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14203_2_lut.init = 16'h2222;
    FD1P3AX read_value__i11 (.D(n30324), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i11.GSR = "ENABLED";
    FD1P3AX read_value__i12 (.D(n30323), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i12.GSR = "ENABLED";
    FD1P3AX read_value__i13 (.D(n30322), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i13.GSR = "ENABLED";
    FD1P3AX read_value__i14 (.D(n30321), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i14.GSR = "ENABLED";
    LUT4 i11580_3_lut (.A(div_factor_reg[4]), .B(steps_reg[4]), .C(\register_addr[0] ), 
         .Z(n2_adj_4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(460[13:26])
    defparam i11580_3_lut.init = 16'hcaca;
    LUT4 i24495_3_lut (.A(Stepper_X_M1_c_1), .B(fault_latched), .C(\register_addr[0] ), 
         .Z(n30854)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24495_3_lut.init = 16'hcaca;
    LUT4 i14202_2_lut (.A(Stepper_X_Dir_c), .B(\register_addr[0] ), .Z(n1_adj_5)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam i14202_2_lut.init = 16'h2222;
    LUT4 i24496_3_lut (.A(div_factor_reg[1]), .B(steps_reg[1]), .C(\register_addr[0] ), 
         .Z(n30855)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24496_3_lut.init = 16'hcaca;
    FD1P3IX read_value__i0 (.D(n30865), .SP(n11966), .CD(n32354), .CK(debug_c_c), 
            .Q(read_value[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i0.GSR = "ENABLED";
    LUT4 mux_1600_Mux_5_i2_3_lut (.A(div_factor_reg[5]), .B(steps_reg[5]), 
         .C(\register_addr[0] ), .Z(n2_adj_6)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(84[8] 110[15])
    defparam mux_1600_Mux_5_i2_3_lut.init = 16'hcaca;
    PFUMX i24494 (.BLUT(n30851), .ALUT(n30852), .C0(\register_addr[1] ), 
          .Z(n30853));
    FD1P3AX read_value__i15 (.D(n30320), .SP(n11966), .CK(debug_c_c), 
            .Q(read_value[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam read_value__i15.GSR = "ENABLED";
    IFS1P3DX fault_latched_178 (.D(Stepper_X_nFault_c), .SP(VCC_net), .SCLK(debug_c_c), 
            .CD(GND_net), .Q(fault_latched)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=25, LSE_RCOL=45, LSE_LLINE=559, LSE_RLINE=572 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam fault_latched_178.GSR = "ENABLED";
    PFUMX i24497 (.BLUT(n30854), .ALUT(n30855), .C0(\register_addr[1] ), 
          .Z(n30856));
    PFUMX mux_1600_Mux_6_i3 (.BLUT(n1), .ALUT(n2), .C0(\register_addr[1] ), 
          .Z(n5188[6]));
    LUT4 i24504_3_lut (.A(Stepper_X_M0_c_0), .B(div_factor_reg[0]), .C(\register_addr[1] ), 
         .Z(n30863)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24504_3_lut.init = 16'hcaca;
    LUT4 i24505_3_lut (.A(n21), .B(steps_reg[0]), .C(\register_addr[1] ), 
         .Z(n30864)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24505_3_lut.init = 16'hcaca;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n28332)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(steps_reg[8]), .B(steps_reg[18]), .C(steps_reg[28]), 
         .D(steps_reg[24]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(steps_reg[26]), .B(n52), .C(n38), .D(steps_reg[9]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(steps_reg[4]), .B(steps_reg[21]), .C(steps_reg[11]), 
         .D(steps_reg[25]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(steps_reg[30]), .B(\steps_reg[7] ), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(steps_reg[0]), .B(n56), .C(n46), .D(steps_reg[1]), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_17 (.A(div_factor_reg[8]), .B(n30313), .C(steps_reg[8]), 
         .D(\register_addr[0] ), .Z(n30327)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_17.init = 16'hc088;
    LUT4 i22_4_lut (.A(steps_reg[22]), .B(steps_reg[6]), .C(steps_reg[5]), 
         .D(steps_reg[10]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(steps_reg[14]), .B(steps_reg[19]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i24_4_lut (.A(steps_reg[29]), .B(steps_reg[3]), .C(steps_reg[13]), 
         .D(steps_reg[31]), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(steps_reg[15]), .B(steps_reg[23]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(steps_reg[16]), .B(steps_reg[20]), .C(steps_reg[2]), 
         .D(steps_reg[27]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut (.A(n32448), .B(n32379), .C(n32504), .D(n30401), .Z(n8048)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_4_lut.init = 16'h0400;
    LUT4 i6_2_lut (.A(steps_reg[12]), .B(steps_reg[17]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    PFUMX i11575 (.BLUT(n17324), .ALUT(n13), .C0(\register_addr[0] ), 
          .Z(n5188[7]));
    LUT4 i1_2_lut_adj_18 (.A(int_step), .B(control_reg[3]), .Z(Stepper_X_Step_c)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut_adj_18.init = 16'h9999;
    LUT4 i1_4_lut_adj_19 (.A(div_factor_reg[9]), .B(n30313), .C(steps_reg[9]), 
         .D(\register_addr[0] ), .Z(n30326)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_19.init = 16'hc088;
    LUT4 i1_4_lut_adj_20 (.A(div_factor_reg[10]), .B(n30313), .C(steps_reg[10]), 
         .D(\register_addr[0] ), .Z(n30325)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_20.init = 16'hc088;
    LUT4 i1_4_lut_adj_21 (.A(div_factor_reg[11]), .B(n30313), .C(steps_reg[11]), 
         .D(\register_addr[0] ), .Z(n30324)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_21.init = 16'hc088;
    LUT4 i1_4_lut_adj_22 (.A(div_factor_reg[12]), .B(n30313), .C(steps_reg[12]), 
         .D(\register_addr[0] ), .Z(n30323)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_22.init = 16'hc088;
    LUT4 i1_4_lut_adj_23 (.A(div_factor_reg[13]), .B(n30313), .C(steps_reg[13]), 
         .D(\register_addr[0] ), .Z(n30322)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_23.init = 16'hc088;
    LUT4 i1_4_lut_adj_24 (.A(div_factor_reg[14]), .B(n30313), .C(steps_reg[14]), 
         .D(\register_addr[0] ), .Z(n30321)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_24.init = 16'hc088;
    LUT4 i24492_3_lut (.A(Stepper_X_M2_c_2), .B(limit_latched), .C(\register_addr[0] ), 
         .Z(n30851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24492_3_lut.init = 16'hcaca;
    LUT4 i24493_3_lut (.A(div_factor_reg[2]), .B(steps_reg[2]), .C(\register_addr[0] ), 
         .Z(n30852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24493_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_25 (.A(div_factor_reg[15]), .B(n30313), .C(steps_reg[15]), 
         .D(\register_addr[0] ), .Z(n30320)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(58[9] 128[6])
    defparam i1_4_lut_adj_25.init = 16'hc088;
    CCU2D sub_125_add_2_33 (.A0(steps_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27757), .S0(n224[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_33.INIT0 = 16'h5555;
    defparam sub_125_add_2_33.INIT1 = 16'h0000;
    defparam sub_125_add_2_33.INJECT1_0 = "NO";
    defparam sub_125_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_31 (.A0(steps_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27756), .COUT(n27757), .S0(n224[29]), 
          .S1(n224[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_31.INIT0 = 16'h5555;
    defparam sub_125_add_2_31.INIT1 = 16'h5555;
    defparam sub_125_add_2_31.INJECT1_0 = "NO";
    defparam sub_125_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_29 (.A0(steps_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27755), .COUT(n27756), .S0(n224[27]), 
          .S1(n224[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_29.INIT0 = 16'h5555;
    defparam sub_125_add_2_29.INIT1 = 16'h5555;
    defparam sub_125_add_2_29.INJECT1_0 = "NO";
    defparam sub_125_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_27 (.A0(steps_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27754), .COUT(n27755), .S0(n224[25]), 
          .S1(n224[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_27.INIT0 = 16'h5555;
    defparam sub_125_add_2_27.INIT1 = 16'h5555;
    defparam sub_125_add_2_27.INJECT1_0 = "NO";
    defparam sub_125_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_25 (.A0(steps_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27753), .COUT(n27754), .S0(n224[23]), 
          .S1(n224[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_25.INIT0 = 16'h5555;
    defparam sub_125_add_2_25.INIT1 = 16'h5555;
    defparam sub_125_add_2_25.INJECT1_0 = "NO";
    defparam sub_125_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_23 (.A0(steps_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27752), .COUT(n27753), .S0(n224[21]), 
          .S1(n224[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_23.INIT0 = 16'h5555;
    defparam sub_125_add_2_23.INIT1 = 16'h5555;
    defparam sub_125_add_2_23.INJECT1_0 = "NO";
    defparam sub_125_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_21 (.A0(steps_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27751), .COUT(n27752), .S0(n224[19]), 
          .S1(n224[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_21.INIT0 = 16'h5555;
    defparam sub_125_add_2_21.INIT1 = 16'h5555;
    defparam sub_125_add_2_21.INJECT1_0 = "NO";
    defparam sub_125_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_19 (.A0(steps_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27750), .COUT(n27751), .S0(n224[17]), 
          .S1(n224[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_19.INIT0 = 16'h5555;
    defparam sub_125_add_2_19.INIT1 = 16'h5555;
    defparam sub_125_add_2_19.INJECT1_0 = "NO";
    defparam sub_125_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_17 (.A0(steps_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27749), .COUT(n27750), .S0(n224[15]), 
          .S1(n224[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_17.INIT0 = 16'h5555;
    defparam sub_125_add_2_17.INIT1 = 16'h5555;
    defparam sub_125_add_2_17.INJECT1_0 = "NO";
    defparam sub_125_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_15 (.A0(steps_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27748), .COUT(n27749), .S0(n224[13]), 
          .S1(n224[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_15.INIT0 = 16'h5555;
    defparam sub_125_add_2_15.INIT1 = 16'h5555;
    defparam sub_125_add_2_15.INJECT1_0 = "NO";
    defparam sub_125_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_125_add_2_13 (.A0(steps_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(steps_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27747), .COUT(n27748), .S0(n224[11]), 
          .S1(n224[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(79[21:34])
    defparam sub_125_add_2_13.INIT0 = 16'h5555;
    defparam sub_125_add_2_13.INIT1 = 16'h5555;
    defparam sub_125_add_2_13.INJECT1_0 = "NO";
    defparam sub_125_add_2_13.INJECT1_1 = "NO";
    ClockDivider_U8 step_clk_gen (.step_clk(step_clk), .debug_c_c(debug_c_c), 
            .n32433(n32433), .n34320(n34320), .prev_step_clk(prev_step_clk), 
            .n21(n21), .n32362(n32362), .n12(n12), .GND_net(GND_net), 
            .div_factor_reg({div_factor_reg})) /* synthesis syn_module_defined=1 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/arm.v(129[15] 132[42])
    
endmodule
//
// Verilog Description of module ClockDivider_U8
//

module ClockDivider_U8 (step_clk, debug_c_c, n32433, n34320, prev_step_clk, 
            n21, n32362, n12, GND_net, div_factor_reg) /* synthesis syn_module_defined=1 */ ;
    output step_clk;
    input debug_c_c;
    input n32433;
    input n34320;
    input prev_step_clk;
    input n21;
    output n32362;
    output n12;
    input GND_net;
    input [31:0]div_factor_reg;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire n6813, n6848, n32337, n6882, n14150;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    wire [31:0]n134;
    
    wire n27693;
    wire [31:0]int_factor;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(45[13:23])
    wire [31:0]n40;
    
    wire n27692, n27691, n27690, n27689, n27688, n27687, n27686, 
        n27685, n27684, n27683, n27682, n27681, n27680, n27679, 
        n27505, n27504, n27678, n27503, n27502, n27501, n27500, 
        n27499, n27498, n27497, n27496, n27495, n27494, n27493, 
        n27492, n27491, n27490, n27489, n27488, n27487, n27486, 
        n27485, n27484, n27483, n27482, n27481, n27480, n27479, 
        n27478, n27477, n27476, n27475, n27474, n27473, n27472, 
        n27471, n27470, n27469, n27468, n27467, n27466, n27465, 
        n27464, n27463, n27462, n27461, n27460, n27459, n27458, 
        n27861, n27860, n27859, n27858, n27857, n27856, n27855, 
        n27854, n27853, n27852, n27851, n27850, n27849, n27848, 
        n27847, n27846;
    
    FD1S3IX clk_o_22 (.D(n6813), .CK(debug_c_c), .CD(n32433), .Q(step_clk));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    LUT4 i954_2_lut_rep_243 (.A(n6848), .B(n34320), .Z(n32337)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i954_2_lut_rep_243.init = 16'heeee;
    LUT4 i8470_2_lut_3_lut (.A(n6848), .B(n34320), .C(n6882), .Z(n14150)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i8470_2_lut_3_lut.init = 16'he0e0;
    FD1S3IX count_2176__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i0.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_268 (.A(prev_step_clk), .B(n21), .C(step_clk), .Z(n32362)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam i2_3_lut_rep_268.init = 16'h4040;
    LUT4 i1_4_lut_4_lut (.A(prev_step_clk), .B(n21), .C(step_clk), .D(n34320), 
         .Z(n12)) /* synthesis lut_function=(!(A (C+(D))+!A (((D)+!C)+!B))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam i1_4_lut_4_lut.init = 16'h004a;
    CCU2D sub_7_add_2_33 (.A0(int_factor[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27693), .S0(n40[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_33.INIT0 = 16'h5555;
    defparam sub_7_add_2_33.INIT1 = 16'h0000;
    defparam sub_7_add_2_33.INJECT1_0 = "NO";
    defparam sub_7_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_31 (.A0(int_factor[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27692), .COUT(n27693), .S0(n40[29]), .S1(n40[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_31.INIT0 = 16'h5555;
    defparam sub_7_add_2_31.INIT1 = 16'h5555;
    defparam sub_7_add_2_31.INJECT1_0 = "NO";
    defparam sub_7_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_29 (.A0(int_factor[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27691), .COUT(n27692), .S0(n40[27]), .S1(n40[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_29.INIT0 = 16'h5555;
    defparam sub_7_add_2_29.INIT1 = 16'h5555;
    defparam sub_7_add_2_29.INJECT1_0 = "NO";
    defparam sub_7_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_27 (.A0(int_factor[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27690), .COUT(n27691), .S0(n40[25]), .S1(n40[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_27.INIT0 = 16'h5555;
    defparam sub_7_add_2_27.INIT1 = 16'h5555;
    defparam sub_7_add_2_27.INJECT1_0 = "NO";
    defparam sub_7_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_25 (.A0(int_factor[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27689), .COUT(n27690), .S0(n40[23]), .S1(n40[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_25.INIT0 = 16'h5555;
    defparam sub_7_add_2_25.INIT1 = 16'h5555;
    defparam sub_7_add_2_25.INJECT1_0 = "NO";
    defparam sub_7_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_23 (.A0(int_factor[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27688), .COUT(n27689), .S0(n40[21]), .S1(n40[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_23.INIT0 = 16'h5555;
    defparam sub_7_add_2_23.INIT1 = 16'h5555;
    defparam sub_7_add_2_23.INJECT1_0 = "NO";
    defparam sub_7_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_21 (.A0(int_factor[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27687), .COUT(n27688), .S0(n40[19]), .S1(n40[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_21.INIT0 = 16'h5555;
    defparam sub_7_add_2_21.INIT1 = 16'h5555;
    defparam sub_7_add_2_21.INJECT1_0 = "NO";
    defparam sub_7_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_19 (.A0(int_factor[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27686), .COUT(n27687), .S0(n40[17]), .S1(n40[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_19.INIT0 = 16'h5555;
    defparam sub_7_add_2_19.INIT1 = 16'h5555;
    defparam sub_7_add_2_19.INJECT1_0 = "NO";
    defparam sub_7_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_17 (.A0(int_factor[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27685), .COUT(n27686), .S0(n40[15]), .S1(n40[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_17.INIT0 = 16'h5555;
    defparam sub_7_add_2_17.INIT1 = 16'h5555;
    defparam sub_7_add_2_17.INJECT1_0 = "NO";
    defparam sub_7_add_2_17.INJECT1_1 = "NO";
    FD1P3JX int_factor_i0_i1 (.D(div_factor_reg[1]), .SP(n32337), .PD(n14150), 
            .CK(debug_c_c), .Q(int_factor[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i1.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i2 (.D(div_factor_reg[2]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i2.GSR = "ENABLED";
    CCU2D sub_7_add_2_15 (.A0(int_factor[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27684), .COUT(n27685), .S0(n40[13]), .S1(n40[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_15.INIT0 = 16'h5555;
    defparam sub_7_add_2_15.INIT1 = 16'h5555;
    defparam sub_7_add_2_15.INJECT1_0 = "NO";
    defparam sub_7_add_2_15.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i3 (.D(div_factor_reg[3]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i3.GSR = "ENABLED";
    CCU2D sub_7_add_2_13 (.A0(int_factor[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27683), .COUT(n27684), .S0(n40[11]), .S1(n40[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_13.INIT0 = 16'h5555;
    defparam sub_7_add_2_13.INIT1 = 16'h5555;
    defparam sub_7_add_2_13.INJECT1_0 = "NO";
    defparam sub_7_add_2_13.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i4 (.D(div_factor_reg[4]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i4.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i5 (.D(div_factor_reg[5]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i5.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i6 (.D(div_factor_reg[6]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i6.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i7 (.D(div_factor_reg[7]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i7.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i8 (.D(div_factor_reg[8]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i8.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i9 (.D(div_factor_reg[9]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i9.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i10 (.D(div_factor_reg[10]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i10.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i11 (.D(div_factor_reg[11]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i11.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i12 (.D(div_factor_reg[12]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i12.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i13 (.D(div_factor_reg[13]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i13.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i14 (.D(div_factor_reg[14]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i14.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i15 (.D(div_factor_reg[15]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i15.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i16 (.D(div_factor_reg[16]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i16.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i17 (.D(div_factor_reg[17]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i17.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i18 (.D(div_factor_reg[18]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i18.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i19 (.D(div_factor_reg[19]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i19.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i0 (.D(div_factor_reg[0]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i0.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i20 (.D(div_factor_reg[20]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i20.GSR = "ENABLED";
    CCU2D sub_7_add_2_11 (.A0(int_factor[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27682), .COUT(n27683), .S0(n40[9]), .S1(n40[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_11.INIT0 = 16'h5555;
    defparam sub_7_add_2_11.INIT1 = 16'h5555;
    defparam sub_7_add_2_11.INJECT1_0 = "NO";
    defparam sub_7_add_2_11.INJECT1_1 = "NO";
    FD1S3IX count_2176__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i1.GSR = "ENABLED";
    FD1S3IX count_2176__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i2.GSR = "ENABLED";
    FD1S3IX count_2176__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i3.GSR = "ENABLED";
    FD1S3IX count_2176__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i4.GSR = "ENABLED";
    FD1S3IX count_2176__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i5.GSR = "ENABLED";
    FD1S3IX count_2176__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i6.GSR = "ENABLED";
    FD1S3IX count_2176__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i7.GSR = "ENABLED";
    FD1S3IX count_2176__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i8.GSR = "ENABLED";
    FD1S3IX count_2176__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i9.GSR = "ENABLED";
    FD1S3IX count_2176__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i10.GSR = "ENABLED";
    FD1S3IX count_2176__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i11.GSR = "ENABLED";
    FD1S3IX count_2176__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i12.GSR = "ENABLED";
    FD1S3IX count_2176__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i13.GSR = "ENABLED";
    FD1S3IX count_2176__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i14.GSR = "ENABLED";
    FD1S3IX count_2176__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i15.GSR = "ENABLED";
    FD1S3IX count_2176__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i16.GSR = "ENABLED";
    FD1S3IX count_2176__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i17.GSR = "ENABLED";
    FD1S3IX count_2176__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i18.GSR = "ENABLED";
    FD1S3IX count_2176__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i19.GSR = "ENABLED";
    FD1S3IX count_2176__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i20.GSR = "ENABLED";
    FD1S3IX count_2176__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i21.GSR = "ENABLED";
    FD1S3IX count_2176__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i22.GSR = "ENABLED";
    FD1S3IX count_2176__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i23.GSR = "ENABLED";
    FD1S3IX count_2176__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i24.GSR = "ENABLED";
    FD1S3IX count_2176__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i25.GSR = "ENABLED";
    FD1S3IX count_2176__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i26.GSR = "ENABLED";
    FD1S3IX count_2176__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i27.GSR = "ENABLED";
    FD1S3IX count_2176__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i28.GSR = "ENABLED";
    FD1S3IX count_2176__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i29.GSR = "ENABLED";
    FD1S3IX count_2176__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i30.GSR = "ENABLED";
    FD1S3IX count_2176__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n32337), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176__i31.GSR = "ENABLED";
    CCU2D sub_7_add_2_9 (.A0(int_factor[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27681), .COUT(n27682), .S0(n40[7]), .S1(n40[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_9.INIT0 = 16'h5555;
    defparam sub_7_add_2_9.INIT1 = 16'h5555;
    defparam sub_7_add_2_9.INJECT1_0 = "NO";
    defparam sub_7_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_7 (.A0(int_factor[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27680), .COUT(n27681), .S0(n40[5]), .S1(n40[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_7.INIT0 = 16'h5555;
    defparam sub_7_add_2_7.INIT1 = 16'h5555;
    defparam sub_7_add_2_7.INJECT1_0 = "NO";
    defparam sub_7_add_2_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i21 (.D(div_factor_reg[21]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i21.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i22 (.D(div_factor_reg[22]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i22.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i23 (.D(div_factor_reg[23]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i23.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i24 (.D(div_factor_reg[24]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i24.GSR = "ENABLED";
    CCU2D sub_7_add_2_5 (.A0(int_factor[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27679), .COUT(n27680), .S0(n40[3]), .S1(n40[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_5.INIT0 = 16'h5555;
    defparam sub_7_add_2_5.INIT1 = 16'h5555;
    defparam sub_7_add_2_5.INJECT1_0 = "NO";
    defparam sub_7_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27505), .S1(n6813));
    defparam sub_1714_add_2_33.INIT0 = 16'h5555;
    defparam sub_1714_add_2_33.INIT1 = 16'h0000;
    defparam sub_1714_add_2_33.INJECT1_0 = "NO";
    defparam sub_1714_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_31 (.A0(count[29]), .B0(int_factor[30]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(int_factor[31]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27504), .COUT(n27505));
    defparam sub_1714_add_2_31.INIT0 = 16'h5999;
    defparam sub_1714_add_2_31.INIT1 = 16'h5999;
    defparam sub_1714_add_2_31.INJECT1_0 = "NO";
    defparam sub_1714_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_3 (.A0(int_factor[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(int_factor[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27678), .COUT(n27679), .S0(n40[1]), .S1(n40[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_3.INIT0 = 16'h5555;
    defparam sub_7_add_2_3.INIT1 = 16'h5555;
    defparam sub_7_add_2_3.INJECT1_0 = "NO";
    defparam sub_7_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_29 (.A0(count[27]), .B0(int_factor[28]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(int_factor[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27503), .COUT(n27504));
    defparam sub_1714_add_2_29.INIT0 = 16'h5999;
    defparam sub_1714_add_2_29.INIT1 = 16'h5999;
    defparam sub_1714_add_2_29.INJECT1_0 = "NO";
    defparam sub_1714_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_7_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(int_factor[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27678), .S1(n40[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(65[18:30])
    defparam sub_7_add_2_1.INIT0 = 16'hF000;
    defparam sub_7_add_2_1.INIT1 = 16'h5555;
    defparam sub_7_add_2_1.INJECT1_0 = "NO";
    defparam sub_7_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_27 (.A0(count[25]), .B0(int_factor[26]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(int_factor[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27502), .COUT(n27503));
    defparam sub_1714_add_2_27.INIT0 = 16'h5999;
    defparam sub_1714_add_2_27.INIT1 = 16'h5999;
    defparam sub_1714_add_2_27.INJECT1_0 = "NO";
    defparam sub_1714_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_25 (.A0(count[23]), .B0(int_factor[24]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(int_factor[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27501), .COUT(n27502));
    defparam sub_1714_add_2_25.INIT0 = 16'h5999;
    defparam sub_1714_add_2_25.INIT1 = 16'h5999;
    defparam sub_1714_add_2_25.INJECT1_0 = "NO";
    defparam sub_1714_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_23 (.A0(count[21]), .B0(int_factor[22]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(int_factor[23]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27500), .COUT(n27501));
    defparam sub_1714_add_2_23.INIT0 = 16'h5999;
    defparam sub_1714_add_2_23.INIT1 = 16'h5999;
    defparam sub_1714_add_2_23.INJECT1_0 = "NO";
    defparam sub_1714_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_21 (.A0(count[19]), .B0(int_factor[20]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(int_factor[21]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27499), .COUT(n27500));
    defparam sub_1714_add_2_21.INIT0 = 16'h5999;
    defparam sub_1714_add_2_21.INIT1 = 16'h5999;
    defparam sub_1714_add_2_21.INJECT1_0 = "NO";
    defparam sub_1714_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_19 (.A0(count[17]), .B0(int_factor[18]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(int_factor[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27498), .COUT(n27499));
    defparam sub_1714_add_2_19.INIT0 = 16'h5999;
    defparam sub_1714_add_2_19.INIT1 = 16'h5999;
    defparam sub_1714_add_2_19.INJECT1_0 = "NO";
    defparam sub_1714_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_17 (.A0(count[15]), .B0(int_factor[16]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(int_factor[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27497), .COUT(n27498));
    defparam sub_1714_add_2_17.INIT0 = 16'h5999;
    defparam sub_1714_add_2_17.INIT1 = 16'h5999;
    defparam sub_1714_add_2_17.INJECT1_0 = "NO";
    defparam sub_1714_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_15 (.A0(count[13]), .B0(int_factor[14]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(int_factor[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27496), .COUT(n27497));
    defparam sub_1714_add_2_15.INIT0 = 16'h5999;
    defparam sub_1714_add_2_15.INIT1 = 16'h5999;
    defparam sub_1714_add_2_15.INJECT1_0 = "NO";
    defparam sub_1714_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_13 (.A0(count[11]), .B0(int_factor[12]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(int_factor[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27495), .COUT(n27496));
    defparam sub_1714_add_2_13.INIT0 = 16'h5999;
    defparam sub_1714_add_2_13.INIT1 = 16'h5999;
    defparam sub_1714_add_2_13.INJECT1_0 = "NO";
    defparam sub_1714_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_11 (.A0(count[9]), .B0(int_factor[10]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(int_factor[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27494), .COUT(n27495));
    defparam sub_1714_add_2_11.INIT0 = 16'h5999;
    defparam sub_1714_add_2_11.INIT1 = 16'h5999;
    defparam sub_1714_add_2_11.INJECT1_0 = "NO";
    defparam sub_1714_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_9 (.A0(count[7]), .B0(int_factor[8]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(int_factor[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27493), .COUT(n27494));
    defparam sub_1714_add_2_9.INIT0 = 16'h5999;
    defparam sub_1714_add_2_9.INIT1 = 16'h5999;
    defparam sub_1714_add_2_9.INJECT1_0 = "NO";
    defparam sub_1714_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_7 (.A0(count[5]), .B0(int_factor[6]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(int_factor[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27492), .COUT(n27493));
    defparam sub_1714_add_2_7.INIT0 = 16'h5999;
    defparam sub_1714_add_2_7.INIT1 = 16'h5999;
    defparam sub_1714_add_2_7.INJECT1_0 = "NO";
    defparam sub_1714_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_5 (.A0(count[3]), .B0(int_factor[4]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(int_factor[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27491), .COUT(n27492));
    defparam sub_1714_add_2_5.INIT0 = 16'h5999;
    defparam sub_1714_add_2_5.INIT1 = 16'h5999;
    defparam sub_1714_add_2_5.INJECT1_0 = "NO";
    defparam sub_1714_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_3 (.A0(count[1]), .B0(int_factor[2]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(int_factor[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27490), .COUT(n27491));
    defparam sub_1714_add_2_3.INIT0 = 16'h5999;
    defparam sub_1714_add_2_3.INIT1 = 16'h5999;
    defparam sub_1714_add_2_3.INJECT1_0 = "NO";
    defparam sub_1714_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1714_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(int_factor[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n27490));
    defparam sub_1714_add_2_1.INIT0 = 16'h0000;
    defparam sub_1714_add_2_1.INIT1 = 16'h5999;
    defparam sub_1714_add_2_1.INJECT1_0 = "NO";
    defparam sub_1714_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_33 (.A0(count[31]), .B0(n40[31]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27489), .S1(n6848));
    defparam sub_1716_add_2_33.INIT0 = 16'h5999;
    defparam sub_1716_add_2_33.INIT1 = 16'h0000;
    defparam sub_1716_add_2_33.INJECT1_0 = "NO";
    defparam sub_1716_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_31 (.A0(count[29]), .B0(n40[29]), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(n40[30]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27488), .COUT(n27489));
    defparam sub_1716_add_2_31.INIT0 = 16'h5999;
    defparam sub_1716_add_2_31.INIT1 = 16'h5999;
    defparam sub_1716_add_2_31.INJECT1_0 = "NO";
    defparam sub_1716_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_29 (.A0(count[27]), .B0(n40[27]), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(n40[28]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27487), .COUT(n27488));
    defparam sub_1716_add_2_29.INIT0 = 16'h5999;
    defparam sub_1716_add_2_29.INIT1 = 16'h5999;
    defparam sub_1716_add_2_29.INJECT1_0 = "NO";
    defparam sub_1716_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_27 (.A0(count[25]), .B0(n40[25]), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(n40[26]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27486), .COUT(n27487));
    defparam sub_1716_add_2_27.INIT0 = 16'h5999;
    defparam sub_1716_add_2_27.INIT1 = 16'h5999;
    defparam sub_1716_add_2_27.INJECT1_0 = "NO";
    defparam sub_1716_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_25 (.A0(count[23]), .B0(n40[23]), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(n40[24]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27485), .COUT(n27486));
    defparam sub_1716_add_2_25.INIT0 = 16'h5999;
    defparam sub_1716_add_2_25.INIT1 = 16'h5999;
    defparam sub_1716_add_2_25.INJECT1_0 = "NO";
    defparam sub_1716_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_23 (.A0(count[21]), .B0(n40[21]), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(n40[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27484), .COUT(n27485));
    defparam sub_1716_add_2_23.INIT0 = 16'h5999;
    defparam sub_1716_add_2_23.INIT1 = 16'h5999;
    defparam sub_1716_add_2_23.INJECT1_0 = "NO";
    defparam sub_1716_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_21 (.A0(count[19]), .B0(n40[19]), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(n40[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27483), .COUT(n27484));
    defparam sub_1716_add_2_21.INIT0 = 16'h5999;
    defparam sub_1716_add_2_21.INIT1 = 16'h5999;
    defparam sub_1716_add_2_21.INJECT1_0 = "NO";
    defparam sub_1716_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_19 (.A0(count[17]), .B0(n40[17]), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(n40[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27482), .COUT(n27483));
    defparam sub_1716_add_2_19.INIT0 = 16'h5999;
    defparam sub_1716_add_2_19.INIT1 = 16'h5999;
    defparam sub_1716_add_2_19.INJECT1_0 = "NO";
    defparam sub_1716_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_17 (.A0(count[15]), .B0(n40[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(n40[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27481), .COUT(n27482));
    defparam sub_1716_add_2_17.INIT0 = 16'h5999;
    defparam sub_1716_add_2_17.INIT1 = 16'h5999;
    defparam sub_1716_add_2_17.INJECT1_0 = "NO";
    defparam sub_1716_add_2_17.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i25 (.D(div_factor_reg[25]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i25.GSR = "ENABLED";
    CCU2D sub_1716_add_2_15 (.A0(count[13]), .B0(n40[13]), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(n40[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27480), .COUT(n27481));
    defparam sub_1716_add_2_15.INIT0 = 16'h5999;
    defparam sub_1716_add_2_15.INIT1 = 16'h5999;
    defparam sub_1716_add_2_15.INJECT1_0 = "NO";
    defparam sub_1716_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_13 (.A0(count[11]), .B0(n40[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(n40[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27479), .COUT(n27480));
    defparam sub_1716_add_2_13.INIT0 = 16'h5999;
    defparam sub_1716_add_2_13.INIT1 = 16'h5999;
    defparam sub_1716_add_2_13.INJECT1_0 = "NO";
    defparam sub_1716_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_11 (.A0(count[9]), .B0(n40[9]), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(n40[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n27478), .COUT(n27479));
    defparam sub_1716_add_2_11.INIT0 = 16'h5999;
    defparam sub_1716_add_2_11.INIT1 = 16'h5999;
    defparam sub_1716_add_2_11.INJECT1_0 = "NO";
    defparam sub_1716_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_9 (.A0(count[7]), .B0(n40[7]), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(n40[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27477), .COUT(n27478));
    defparam sub_1716_add_2_9.INIT0 = 16'h5999;
    defparam sub_1716_add_2_9.INIT1 = 16'h5999;
    defparam sub_1716_add_2_9.INJECT1_0 = "NO";
    defparam sub_1716_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_7 (.A0(count[5]), .B0(n40[5]), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(n40[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27476), .COUT(n27477));
    defparam sub_1716_add_2_7.INIT0 = 16'h5999;
    defparam sub_1716_add_2_7.INIT1 = 16'h5999;
    defparam sub_1716_add_2_7.INJECT1_0 = "NO";
    defparam sub_1716_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_5 (.A0(count[3]), .B0(n40[3]), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(n40[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27475), .COUT(n27476));
    defparam sub_1716_add_2_5.INIT0 = 16'h5999;
    defparam sub_1716_add_2_5.INIT1 = 16'h5999;
    defparam sub_1716_add_2_5.INJECT1_0 = "NO";
    defparam sub_1716_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_3 (.A0(count[1]), .B0(n40[1]), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(n40[2]), .C1(GND_net), .D1(GND_net), 
          .CIN(n27474), .COUT(n27475));
    defparam sub_1716_add_2_3.INIT0 = 16'h5999;
    defparam sub_1716_add_2_3.INIT1 = 16'h5999;
    defparam sub_1716_add_2_3.INJECT1_0 = "NO";
    defparam sub_1716_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1716_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(n40[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n27474));
    defparam sub_1716_add_2_1.INIT0 = 16'h0000;
    defparam sub_1716_add_2_1.INIT1 = 16'h5999;
    defparam sub_1716_add_2_1.INJECT1_0 = "NO";
    defparam sub_1716_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_33 (.A0(div_factor_reg[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27473), .S1(n6882));
    defparam sub_1717_add_2_33.INIT0 = 16'hf555;
    defparam sub_1717_add_2_33.INIT1 = 16'h0000;
    defparam sub_1717_add_2_33.INJECT1_0 = "NO";
    defparam sub_1717_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_31 (.A0(div_factor_reg[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27472), .COUT(n27473));
    defparam sub_1717_add_2_31.INIT0 = 16'hf555;
    defparam sub_1717_add_2_31.INIT1 = 16'hf555;
    defparam sub_1717_add_2_31.INJECT1_0 = "NO";
    defparam sub_1717_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_29 (.A0(div_factor_reg[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27471), .COUT(n27472));
    defparam sub_1717_add_2_29.INIT0 = 16'hf555;
    defparam sub_1717_add_2_29.INIT1 = 16'hf555;
    defparam sub_1717_add_2_29.INJECT1_0 = "NO";
    defparam sub_1717_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_27 (.A0(div_factor_reg[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27470), .COUT(n27471));
    defparam sub_1717_add_2_27.INIT0 = 16'hf555;
    defparam sub_1717_add_2_27.INIT1 = 16'hf555;
    defparam sub_1717_add_2_27.INJECT1_0 = "NO";
    defparam sub_1717_add_2_27.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i26 (.D(div_factor_reg[26]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i26.GSR = "ENABLED";
    CCU2D sub_1717_add_2_25 (.A0(div_factor_reg[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27469), .COUT(n27470));
    defparam sub_1717_add_2_25.INIT0 = 16'hf555;
    defparam sub_1717_add_2_25.INIT1 = 16'hf555;
    defparam sub_1717_add_2_25.INJECT1_0 = "NO";
    defparam sub_1717_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_23 (.A0(div_factor_reg[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27468), .COUT(n27469));
    defparam sub_1717_add_2_23.INIT0 = 16'hf555;
    defparam sub_1717_add_2_23.INIT1 = 16'hf555;
    defparam sub_1717_add_2_23.INJECT1_0 = "NO";
    defparam sub_1717_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_21 (.A0(div_factor_reg[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27467), .COUT(n27468));
    defparam sub_1717_add_2_21.INIT0 = 16'hf555;
    defparam sub_1717_add_2_21.INIT1 = 16'hf555;
    defparam sub_1717_add_2_21.INJECT1_0 = "NO";
    defparam sub_1717_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_19 (.A0(div_factor_reg[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27466), .COUT(n27467));
    defparam sub_1717_add_2_19.INIT0 = 16'hf555;
    defparam sub_1717_add_2_19.INIT1 = 16'hf555;
    defparam sub_1717_add_2_19.INJECT1_0 = "NO";
    defparam sub_1717_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_17 (.A0(div_factor_reg[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27465), .COUT(n27466));
    defparam sub_1717_add_2_17.INIT0 = 16'hf555;
    defparam sub_1717_add_2_17.INIT1 = 16'hf555;
    defparam sub_1717_add_2_17.INJECT1_0 = "NO";
    defparam sub_1717_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_15 (.A0(div_factor_reg[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27464), .COUT(n27465));
    defparam sub_1717_add_2_15.INIT0 = 16'hf555;
    defparam sub_1717_add_2_15.INIT1 = 16'hf555;
    defparam sub_1717_add_2_15.INJECT1_0 = "NO";
    defparam sub_1717_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_13 (.A0(div_factor_reg[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27463), .COUT(n27464));
    defparam sub_1717_add_2_13.INIT0 = 16'hf555;
    defparam sub_1717_add_2_13.INIT1 = 16'hf555;
    defparam sub_1717_add_2_13.INJECT1_0 = "NO";
    defparam sub_1717_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_11 (.A0(div_factor_reg[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27462), .COUT(n27463));
    defparam sub_1717_add_2_11.INIT0 = 16'hf555;
    defparam sub_1717_add_2_11.INIT1 = 16'hf555;
    defparam sub_1717_add_2_11.INJECT1_0 = "NO";
    defparam sub_1717_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_9 (.A0(div_factor_reg[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27461), .COUT(n27462));
    defparam sub_1717_add_2_9.INIT0 = 16'hf555;
    defparam sub_1717_add_2_9.INIT1 = 16'hf555;
    defparam sub_1717_add_2_9.INJECT1_0 = "NO";
    defparam sub_1717_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_7 (.A0(div_factor_reg[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27460), .COUT(n27461));
    defparam sub_1717_add_2_7.INIT0 = 16'hf555;
    defparam sub_1717_add_2_7.INIT1 = 16'hf555;
    defparam sub_1717_add_2_7.INJECT1_0 = "NO";
    defparam sub_1717_add_2_7.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i27 (.D(div_factor_reg[27]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i27.GSR = "ENABLED";
    CCU2D sub_1717_add_2_5 (.A0(div_factor_reg[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27459), .COUT(n27460));
    defparam sub_1717_add_2_5.INIT0 = 16'hf555;
    defparam sub_1717_add_2_5.INIT1 = 16'hf555;
    defparam sub_1717_add_2_5.INJECT1_0 = "NO";
    defparam sub_1717_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_3 (.A0(div_factor_reg[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27458), .COUT(n27459));
    defparam sub_1717_add_2_3.INIT0 = 16'hf555;
    defparam sub_1717_add_2_3.INIT1 = 16'hf555;
    defparam sub_1717_add_2_3.INJECT1_0 = "NO";
    defparam sub_1717_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1717_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(div_factor_reg[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n27458));
    defparam sub_1717_add_2_1.INIT0 = 16'h0000;
    defparam sub_1717_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_1717_add_2_1.INJECT1_0 = "NO";
    defparam sub_1717_add_2_1.INJECT1_1 = "NO";
    FD1P3IX int_factor_i0_i28 (.D(div_factor_reg[28]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i28.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i29 (.D(div_factor_reg[29]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i29.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i30 (.D(div_factor_reg[30]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i30.GSR = "ENABLED";
    FD1P3IX int_factor_i0_i31 (.D(div_factor_reg[31]), .SP(n32337), .CD(n14150), 
            .CK(debug_c_c), .Q(int_factor[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=15, LSE_RCOL=42, LSE_LLINE=129, LSE_RLINE=132 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam int_factor_i0_i31.GSR = "ENABLED";
    CCU2D count_2176_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27861), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_33.INIT1 = 16'h0000;
    defparam count_2176_add_4_33.INJECT1_0 = "NO";
    defparam count_2176_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27860), .COUT(n27861), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_31.INJECT1_0 = "NO";
    defparam count_2176_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27859), .COUT(n27860), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_29.INJECT1_0 = "NO";
    defparam count_2176_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27858), .COUT(n27859), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_27.INJECT1_0 = "NO";
    defparam count_2176_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27857), .COUT(n27858), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_25.INJECT1_0 = "NO";
    defparam count_2176_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27856), .COUT(n27857), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_23.INJECT1_0 = "NO";
    defparam count_2176_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27855), .COUT(n27856), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_21.INJECT1_0 = "NO";
    defparam count_2176_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27854), .COUT(n27855), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_19.INJECT1_0 = "NO";
    defparam count_2176_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27853), .COUT(n27854), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_17.INJECT1_0 = "NO";
    defparam count_2176_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27852), .COUT(n27853), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_15.INJECT1_0 = "NO";
    defparam count_2176_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27851), .COUT(n27852), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_13.INJECT1_0 = "NO";
    defparam count_2176_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27850), .COUT(n27851), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_11.INJECT1_0 = "NO";
    defparam count_2176_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27849), .COUT(n27850), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_9.INJECT1_0 = "NO";
    defparam count_2176_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27848), .COUT(n27849), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_7.INJECT1_0 = "NO";
    defparam count_2176_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27847), .COUT(n27848), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_5.INJECT1_0 = "NO";
    defparam count_2176_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27846), .COUT(n27847), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2176_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2176_add_4_3.INJECT1_0 = "NO";
    defparam count_2176_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2176_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27846), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2176_add_4_1.INIT0 = 16'hF000;
    defparam count_2176_add_4_1.INIT1 = 16'h0555;
    defparam count_2176_add_4_1.INJECT1_0 = "NO";
    defparam count_2176_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module ClockDivider_U10
//

module ClockDivider_U10 (debug_c_c, n241, n34320, n6674, n32341, n30913, 
            n12030, n30995, n12031, n30929, n28304, n30911, n28312, 
            n31000, n28317, n31005, n28308, n31024, n28324, n988, 
            n6, n31049, n12841, n30969, n12138, GND_net) /* synthesis syn_module_defined=1 */ ;
    input debug_c_c;
    input n241;
    input n34320;
    output n6674;
    output n32341;
    input n30913;
    output n12030;
    input n30995;
    output n12031;
    input n30929;
    output n28304;
    input n30911;
    output n28312;
    input n31000;
    output n28317;
    input n31005;
    output n28308;
    input n31024;
    output n28324;
    input n988;
    output n6;
    input n31049;
    output n12841;
    input n30969;
    output n12138;
    input GND_net;
    
    wire debug_c_c /* synthesis SET_AS_NETWORK=debug_c_c */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/uniboard.v(367[13:22])
    
    wire clk_255kHz;
    wire [31:0]count;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(44[13:18])
    
    wire n2550;
    wire [31:0]n134;
    
    wire n6709, n27938, n27937, n27936, n27935, n27934, n27933, 
        n27932, n27931, n27930, n27929, n27928, n27927, n27926, 
        n27925, n27924, n27553, n27552, n27551, n27550, n27549, 
        n27548, n27547, n27546, n27545, n27544, n27543, n27542, 
        n27541, n27540, n27539, n27538, n27797, n27796, n27795, 
        n27794, n27793, n27792, n27791, n27790, n27789, n27788, 
        n27787, n27786, n27785, n27784, n27783, n27782;
    
    FD1S3AX clk_o_22 (.D(n241), .CK(debug_c_c), .Q(clk_255kHz)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=15, LSE_RCOL=41, LSE_LLINE=508, LSE_RLINE=511 */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(47[9] 76[6])
    defparam clk_o_22.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_247 (.A(n34320), .B(clk_255kHz), .C(n6674), .Z(n32341)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i2_3_lut_rep_247.init = 16'h1010;
    LUT4 i24646_2_lut_4_lut (.A(n34320), .B(clk_255kHz), .C(n6674), .D(n30913), 
         .Z(n12030)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24646_2_lut_4_lut.init = 16'h1000;
    LUT4 i24728_2_lut_4_lut (.A(n34320), .B(clk_255kHz), .C(n6674), .D(n30995), 
         .Z(n12031)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24728_2_lut_4_lut.init = 16'h1000;
    LUT4 i24662_2_lut_4_lut (.A(n34320), .B(clk_255kHz), .C(n6674), .D(n30929), 
         .Z(n28304)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24662_2_lut_4_lut.init = 16'h1000;
    LUT4 i24644_2_lut_4_lut (.A(n34320), .B(clk_255kHz), .C(n6674), .D(n30911), 
         .Z(n28312)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24644_2_lut_4_lut.init = 16'h1000;
    LUT4 i24733_2_lut_4_lut (.A(n34320), .B(clk_255kHz), .C(n6674), .D(n31000), 
         .Z(n28317)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24733_2_lut_4_lut.init = 16'h1000;
    LUT4 i24738_2_lut_4_lut (.A(n34320), .B(clk_255kHz), .C(n6674), .D(n31005), 
         .Z(n28308)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24738_2_lut_4_lut.init = 16'h1000;
    LUT4 i24757_2_lut_4_lut (.A(n34320), .B(clk_255kHz), .C(n6674), .D(n31024), 
         .Z(n28324)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24757_2_lut_4_lut.init = 16'h1000;
    LUT4 i2_2_lut_4_lut (.A(n34320), .B(clk_255kHz), .C(n6674), .D(n988), 
         .Z(n6)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i2_2_lut_4_lut.init = 16'h1000;
    LUT4 i24782_2_lut_4_lut (.A(n34320), .B(clk_255kHz), .C(n6674), .D(n31049), 
         .Z(n12841)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24782_2_lut_4_lut.init = 16'h1000;
    LUT4 i24702_2_lut_4_lut (.A(n34320), .B(clk_255kHz), .C(n6674), .D(n30969), 
         .Z(n12138)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i24702_2_lut_4_lut.init = 16'h1000;
    FD1S3IX count_2174__i0 (.D(n134[0]), .CK(debug_c_c), .CD(n2550), .Q(count[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i0.GSR = "ENABLED";
    FD1S3IX count_2174__i1 (.D(n134[1]), .CK(debug_c_c), .CD(n2550), .Q(count[1]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i1.GSR = "ENABLED";
    FD1S3IX count_2174__i2 (.D(n134[2]), .CK(debug_c_c), .CD(n2550), .Q(count[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i2.GSR = "ENABLED";
    FD1S3IX count_2174__i3 (.D(n134[3]), .CK(debug_c_c), .CD(n2550), .Q(count[3]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i3.GSR = "ENABLED";
    FD1S3IX count_2174__i4 (.D(n134[4]), .CK(debug_c_c), .CD(n2550), .Q(count[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i4.GSR = "ENABLED";
    FD1S3IX count_2174__i5 (.D(n134[5]), .CK(debug_c_c), .CD(n2550), .Q(count[5]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i5.GSR = "ENABLED";
    FD1S3IX count_2174__i6 (.D(n134[6]), .CK(debug_c_c), .CD(n2550), .Q(count[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i6.GSR = "ENABLED";
    FD1S3IX count_2174__i7 (.D(n134[7]), .CK(debug_c_c), .CD(n2550), .Q(count[7]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i7.GSR = "ENABLED";
    FD1S3IX count_2174__i8 (.D(n134[8]), .CK(debug_c_c), .CD(n2550), .Q(count[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i8.GSR = "ENABLED";
    FD1S3IX count_2174__i9 (.D(n134[9]), .CK(debug_c_c), .CD(n2550), .Q(count[9]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i9.GSR = "ENABLED";
    FD1S3IX count_2174__i10 (.D(n134[10]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i10.GSR = "ENABLED";
    FD1S3IX count_2174__i11 (.D(n134[11]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[11]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i11.GSR = "ENABLED";
    FD1S3IX count_2174__i12 (.D(n134[12]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i12.GSR = "ENABLED";
    FD1S3IX count_2174__i13 (.D(n134[13]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[13]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i13.GSR = "ENABLED";
    FD1S3IX count_2174__i14 (.D(n134[14]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i14.GSR = "ENABLED";
    FD1S3IX count_2174__i15 (.D(n134[15]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[15]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i15.GSR = "ENABLED";
    FD1S3IX count_2174__i16 (.D(n134[16]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i16.GSR = "ENABLED";
    FD1S3IX count_2174__i17 (.D(n134[17]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[17]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i17.GSR = "ENABLED";
    FD1S3IX count_2174__i18 (.D(n134[18]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i18.GSR = "ENABLED";
    FD1S3IX count_2174__i19 (.D(n134[19]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[19]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i19.GSR = "ENABLED";
    FD1S3IX count_2174__i20 (.D(n134[20]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i20.GSR = "ENABLED";
    FD1S3IX count_2174__i21 (.D(n134[21]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[21]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i21.GSR = "ENABLED";
    FD1S3IX count_2174__i22 (.D(n134[22]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i22.GSR = "ENABLED";
    FD1S3IX count_2174__i23 (.D(n134[23]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[23]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i23.GSR = "ENABLED";
    FD1S3IX count_2174__i24 (.D(n134[24]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i24.GSR = "ENABLED";
    FD1S3IX count_2174__i25 (.D(n134[25]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[25]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i25.GSR = "ENABLED";
    FD1S3IX count_2174__i26 (.D(n134[26]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i26.GSR = "ENABLED";
    FD1S3IX count_2174__i27 (.D(n134[27]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[27]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i27.GSR = "ENABLED";
    FD1S3IX count_2174__i28 (.D(n134[28]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i28.GSR = "ENABLED";
    FD1S3IX count_2174__i29 (.D(n134[29]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[29]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i29.GSR = "ENABLED";
    FD1S3IX count_2174__i30 (.D(n134[30]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i30.GSR = "ENABLED";
    FD1S3IX count_2174__i31 (.D(n134[31]), .CK(debug_c_c), .CD(n2550), 
            .Q(count[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174__i31.GSR = "ENABLED";
    LUT4 i893_2_lut (.A(n6709), .B(n34320), .Z(n2550)) /* synthesis lut_function=(A+(B)) */ ;   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(59[5] 75[8])
    defparam i893_2_lut.init = 16'heeee;
    CCU2D add_21584_32 (.A0(count[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27938), 
          .S1(n6674));
    defparam add_21584_32.INIT0 = 16'h5555;
    defparam add_21584_32.INIT1 = 16'h0000;
    defparam add_21584_32.INJECT1_0 = "NO";
    defparam add_21584_32.INJECT1_1 = "NO";
    CCU2D add_21584_30 (.A0(count[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27937), .COUT(n27938));
    defparam add_21584_30.INIT0 = 16'h5555;
    defparam add_21584_30.INIT1 = 16'h5555;
    defparam add_21584_30.INJECT1_0 = "NO";
    defparam add_21584_30.INJECT1_1 = "NO";
    CCU2D add_21584_28 (.A0(count[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27936), .COUT(n27937));
    defparam add_21584_28.INIT0 = 16'h5555;
    defparam add_21584_28.INIT1 = 16'h5555;
    defparam add_21584_28.INJECT1_0 = "NO";
    defparam add_21584_28.INJECT1_1 = "NO";
    CCU2D add_21584_26 (.A0(count[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27935), .COUT(n27936));
    defparam add_21584_26.INIT0 = 16'h5555;
    defparam add_21584_26.INIT1 = 16'h5555;
    defparam add_21584_26.INJECT1_0 = "NO";
    defparam add_21584_26.INJECT1_1 = "NO";
    CCU2D add_21584_24 (.A0(count[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27934), .COUT(n27935));
    defparam add_21584_24.INIT0 = 16'h5555;
    defparam add_21584_24.INIT1 = 16'h5555;
    defparam add_21584_24.INJECT1_0 = "NO";
    defparam add_21584_24.INJECT1_1 = "NO";
    CCU2D add_21584_22 (.A0(count[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27933), .COUT(n27934));
    defparam add_21584_22.INIT0 = 16'h5555;
    defparam add_21584_22.INIT1 = 16'h5555;
    defparam add_21584_22.INJECT1_0 = "NO";
    defparam add_21584_22.INJECT1_1 = "NO";
    CCU2D add_21584_20 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27932), .COUT(n27933));
    defparam add_21584_20.INIT0 = 16'h5555;
    defparam add_21584_20.INIT1 = 16'h5555;
    defparam add_21584_20.INJECT1_0 = "NO";
    defparam add_21584_20.INJECT1_1 = "NO";
    CCU2D add_21584_18 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27931), .COUT(n27932));
    defparam add_21584_18.INIT0 = 16'h5555;
    defparam add_21584_18.INIT1 = 16'h5555;
    defparam add_21584_18.INJECT1_0 = "NO";
    defparam add_21584_18.INJECT1_1 = "NO";
    CCU2D add_21584_16 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27930), .COUT(n27931));
    defparam add_21584_16.INIT0 = 16'h5555;
    defparam add_21584_16.INIT1 = 16'h5555;
    defparam add_21584_16.INJECT1_0 = "NO";
    defparam add_21584_16.INJECT1_1 = "NO";
    CCU2D add_21584_14 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27929), .COUT(n27930));
    defparam add_21584_14.INIT0 = 16'h5555;
    defparam add_21584_14.INIT1 = 16'h5555;
    defparam add_21584_14.INJECT1_0 = "NO";
    defparam add_21584_14.INJECT1_1 = "NO";
    CCU2D add_21584_12 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27928), .COUT(n27929));
    defparam add_21584_12.INIT0 = 16'h5555;
    defparam add_21584_12.INIT1 = 16'h5555;
    defparam add_21584_12.INJECT1_0 = "NO";
    defparam add_21584_12.INJECT1_1 = "NO";
    CCU2D add_21584_10 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27927), .COUT(n27928));
    defparam add_21584_10.INIT0 = 16'h5555;
    defparam add_21584_10.INIT1 = 16'h5555;
    defparam add_21584_10.INJECT1_0 = "NO";
    defparam add_21584_10.INJECT1_1 = "NO";
    CCU2D add_21584_8 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27926), 
          .COUT(n27927));
    defparam add_21584_8.INIT0 = 16'h5555;
    defparam add_21584_8.INIT1 = 16'h5555;
    defparam add_21584_8.INJECT1_0 = "NO";
    defparam add_21584_8.INJECT1_1 = "NO";
    CCU2D add_21584_6 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27925), 
          .COUT(n27926));
    defparam add_21584_6.INIT0 = 16'h5555;
    defparam add_21584_6.INIT1 = 16'h5555;
    defparam add_21584_6.INJECT1_0 = "NO";
    defparam add_21584_6.INJECT1_1 = "NO";
    CCU2D add_21584_4 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27924), 
          .COUT(n27925));
    defparam add_21584_4.INIT0 = 16'h5555;
    defparam add_21584_4.INIT1 = 16'h5aaa;
    defparam add_21584_4.INJECT1_0 = "NO";
    defparam add_21584_4.INJECT1_1 = "NO";
    CCU2D add_21584_2 (.A0(count[1]), .B0(count[0]), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n27924));
    defparam add_21584_2.INIT0 = 16'h7000;
    defparam add_21584_2.INIT1 = 16'h5aaa;
    defparam add_21584_2.INJECT1_0 = "NO";
    defparam add_21584_2.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27553), .S0(n6709));
    defparam sub_1709_add_2_cout.INIT0 = 16'h0000;
    defparam sub_1709_add_2_cout.INIT1 = 16'h0000;
    defparam sub_1709_add_2_cout.INJECT1_0 = "NO";
    defparam sub_1709_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_32 (.A0(count[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27552), .COUT(n27553));
    defparam sub_1709_add_2_32.INIT0 = 16'h5555;
    defparam sub_1709_add_2_32.INIT1 = 16'h5555;
    defparam sub_1709_add_2_32.INJECT1_0 = "NO";
    defparam sub_1709_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_30 (.A0(count[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27551), .COUT(n27552));
    defparam sub_1709_add_2_30.INIT0 = 16'h5555;
    defparam sub_1709_add_2_30.INIT1 = 16'h5555;
    defparam sub_1709_add_2_30.INJECT1_0 = "NO";
    defparam sub_1709_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_28 (.A0(count[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27550), .COUT(n27551));
    defparam sub_1709_add_2_28.INIT0 = 16'h5555;
    defparam sub_1709_add_2_28.INIT1 = 16'h5555;
    defparam sub_1709_add_2_28.INJECT1_0 = "NO";
    defparam sub_1709_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_26 (.A0(count[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27549), .COUT(n27550));
    defparam sub_1709_add_2_26.INIT0 = 16'h5555;
    defparam sub_1709_add_2_26.INIT1 = 16'h5555;
    defparam sub_1709_add_2_26.INJECT1_0 = "NO";
    defparam sub_1709_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_24 (.A0(count[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27548), .COUT(n27549));
    defparam sub_1709_add_2_24.INIT0 = 16'h5555;
    defparam sub_1709_add_2_24.INIT1 = 16'h5555;
    defparam sub_1709_add_2_24.INJECT1_0 = "NO";
    defparam sub_1709_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_22 (.A0(count[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27547), .COUT(n27548));
    defparam sub_1709_add_2_22.INIT0 = 16'h5555;
    defparam sub_1709_add_2_22.INIT1 = 16'h5555;
    defparam sub_1709_add_2_22.INJECT1_0 = "NO";
    defparam sub_1709_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_20 (.A0(count[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27546), .COUT(n27547));
    defparam sub_1709_add_2_20.INIT0 = 16'h5555;
    defparam sub_1709_add_2_20.INIT1 = 16'h5555;
    defparam sub_1709_add_2_20.INJECT1_0 = "NO";
    defparam sub_1709_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_18 (.A0(count[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27545), .COUT(n27546));
    defparam sub_1709_add_2_18.INIT0 = 16'h5555;
    defparam sub_1709_add_2_18.INIT1 = 16'h5555;
    defparam sub_1709_add_2_18.INJECT1_0 = "NO";
    defparam sub_1709_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_16 (.A0(count[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27544), .COUT(n27545));
    defparam sub_1709_add_2_16.INIT0 = 16'h5555;
    defparam sub_1709_add_2_16.INIT1 = 16'h5555;
    defparam sub_1709_add_2_16.INJECT1_0 = "NO";
    defparam sub_1709_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_14 (.A0(count[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27543), .COUT(n27544));
    defparam sub_1709_add_2_14.INIT0 = 16'h5555;
    defparam sub_1709_add_2_14.INIT1 = 16'h5555;
    defparam sub_1709_add_2_14.INJECT1_0 = "NO";
    defparam sub_1709_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_12 (.A0(count[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27542), .COUT(n27543));
    defparam sub_1709_add_2_12.INIT0 = 16'h5555;
    defparam sub_1709_add_2_12.INIT1 = 16'h5555;
    defparam sub_1709_add_2_12.INJECT1_0 = "NO";
    defparam sub_1709_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_10 (.A0(count[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27541), .COUT(n27542));
    defparam sub_1709_add_2_10.INIT0 = 16'h5555;
    defparam sub_1709_add_2_10.INIT1 = 16'h5555;
    defparam sub_1709_add_2_10.INJECT1_0 = "NO";
    defparam sub_1709_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_8 (.A0(count[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27540), .COUT(n27541));
    defparam sub_1709_add_2_8.INIT0 = 16'h5555;
    defparam sub_1709_add_2_8.INIT1 = 16'h5555;
    defparam sub_1709_add_2_8.INJECT1_0 = "NO";
    defparam sub_1709_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_6 (.A0(count[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27539), .COUT(n27540));
    defparam sub_1709_add_2_6.INIT0 = 16'h5555;
    defparam sub_1709_add_2_6.INIT1 = 16'h5aaa;
    defparam sub_1709_add_2_6.INJECT1_0 = "NO";
    defparam sub_1709_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_4 (.A0(count[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27538), .COUT(n27539));
    defparam sub_1709_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_1709_add_2_4.INIT1 = 16'h5aaa;
    defparam sub_1709_add_2_4.INJECT1_0 = "NO";
    defparam sub_1709_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_1709_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27538));
    defparam sub_1709_add_2_2.INIT0 = 16'h0000;
    defparam sub_1709_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_1709_add_2_2.INJECT1_0 = "NO";
    defparam sub_1709_add_2_2.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_33 (.A0(count[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27797), .S0(n134[31]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_33.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_33.INIT1 = 16'h0000;
    defparam count_2174_add_4_33.INJECT1_0 = "NO";
    defparam count_2174_add_4_33.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_31 (.A0(count[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27796), .COUT(n27797), .S0(n134[29]), 
          .S1(n134[30]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_31.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_31.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_31.INJECT1_0 = "NO";
    defparam count_2174_add_4_31.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_29 (.A0(count[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27795), .COUT(n27796), .S0(n134[27]), 
          .S1(n134[28]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_29.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_29.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_29.INJECT1_0 = "NO";
    defparam count_2174_add_4_29.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_27 (.A0(count[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27794), .COUT(n27795), .S0(n134[25]), 
          .S1(n134[26]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_27.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_27.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_27.INJECT1_0 = "NO";
    defparam count_2174_add_4_27.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_25 (.A0(count[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27793), .COUT(n27794), .S0(n134[23]), 
          .S1(n134[24]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_25.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_25.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_25.INJECT1_0 = "NO";
    defparam count_2174_add_4_25.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_23 (.A0(count[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27792), .COUT(n27793), .S0(n134[21]), 
          .S1(n134[22]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_23.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_23.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_23.INJECT1_0 = "NO";
    defparam count_2174_add_4_23.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27791), .COUT(n27792), .S0(n134[19]), 
          .S1(n134[20]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_21.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_21.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_21.INJECT1_0 = "NO";
    defparam count_2174_add_4_21.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27790), .COUT(n27791), .S0(n134[17]), 
          .S1(n134[18]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_19.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_19.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_19.INJECT1_0 = "NO";
    defparam count_2174_add_4_19.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27789), .COUT(n27790), .S0(n134[15]), 
          .S1(n134[16]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_17.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_17.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_17.INJECT1_0 = "NO";
    defparam count_2174_add_4_17.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27788), .COUT(n27789), .S0(n134[13]), 
          .S1(n134[14]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_15.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_15.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_15.INJECT1_0 = "NO";
    defparam count_2174_add_4_15.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27787), .COUT(n27788), .S0(n134[11]), 
          .S1(n134[12]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_13.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_13.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_13.INJECT1_0 = "NO";
    defparam count_2174_add_4_13.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n27786), .COUT(n27787), .S0(n134[9]), .S1(n134[10]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_11.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_11.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_11.INJECT1_0 = "NO";
    defparam count_2174_add_4_11.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27785), .COUT(n27786), .S0(n134[7]), .S1(n134[8]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_9.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_9.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_9.INJECT1_0 = "NO";
    defparam count_2174_add_4_9.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27784), .COUT(n27785), .S0(n134[5]), .S1(n134[6]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_7.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_7.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_7.INJECT1_0 = "NO";
    defparam count_2174_add_4_7.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27783), .COUT(n27784), .S0(n134[3]), .S1(n134[4]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_5.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_5.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_5.INJECT1_0 = "NO";
    defparam count_2174_add_4_5.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27782), .COUT(n27783), .S0(n134[1]), .S1(n134[2]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_3.INIT0 = 16'hfaaa;
    defparam count_2174_add_4_3.INIT1 = 16'hfaaa;
    defparam count_2174_add_4_3.INJECT1_0 = "NO";
    defparam count_2174_add_4_3.INJECT1_1 = "NO";
    CCU2D count_2174_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n27782), .S1(n134[0]));   // /home/nick/Desktop/nickfolder/documents/projects/in-progress/project 5l - OSURC Rover 2016/electrical/uniboard/software/hdl-verilog/clk.v(74[16:25])
    defparam count_2174_add_4_1.INIT0 = 16'hF000;
    defparam count_2174_add_4_1.INIT1 = 16'h0555;
    defparam count_2174_add_4_1.INJECT1_0 = "NO";
    defparam count_2174_add_4_1.INJECT1_1 = "NO";
    
endmodule
